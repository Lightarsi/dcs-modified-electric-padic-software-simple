*** SPICE deck for cell 5400TP094NEW{sch} from library 5400TP094
*** Created on Сб мар 24, 2018 14:37:07
*** Last revised on Пн сен 10, 2018 14:41:19
*** Written on Пн сен 10, 2018 15:00:08 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
.options parhier=local

*** SUBCIRCUIT basic__key FROM CELL basic:key{sch}
.SUBCKT basic__key M1 M2 X Y adr=0
** GLOBAL gnd
Rres@4 gnd M2 100k
*
*
*
*
Xswitch_m@2 X Y M2 switch_man
.SUBCKT switch_man X Y man
S1 X Y man 0 switch1 OFF
.model switch1 sw vt=2.5 vh=1 ron=500 roff=1000G
.ENDS switch_man
******************************************************
Vvsource@0 M1 0 5

* Spice Code nodes in cell cell 'basic:key{sch}'
.param adr = 67
.ENDS basic__key

*** SUBCIRCUIT _5400TP094__CB FROM CELL CB{sch}
.SUBCKT _5400TP094__CB K0 K1 K10 K11 K12 K13 K2 K3 K4 K5 K6 K7 K8 K9 mAd000_1 mAd000_2 mAd001_1 mAd001_2 mAd002_1 mAd002_2 mAd003_1 mAd003_2 mAd004_1 mAd004_2 mAd005_1 mAd005_2 mAd006_1 mAd006_2 mAd007_1 mAd007_2 mAd010_1 mAd010_2 mAd011_1 mAd011_2 mAd012_1 mAd012_2 mAd013_1 mAd013_2 mAd014_1 mAd014_2 mAd015_1 mAd015_2 mAd016_1 mAd016_2 mAd017_1 mAd017_2 mAd020_1 mAd020_2 mAd021_1 mAd021_2 mAd022_1 mAd022_2 mAd023_1 mAd023_2 mAd024_1 mAd024_2 mAd025_1 mAd025_2 mAd026_1 mAd026_2 mAd027_1 mAd027_2 mAd030_1 
+mAd030_2 mAd031_1 mAd031_2 mAd032_1 mAd032_2 mAd033_1 mAd033_2 mAd034_1 mAd034_2 mAd035_1 mAd035_2 mAd036_1 mAd036_2 mAd037_1 mAd037_2 mAd040_1 mAd040_2 mAd041_1 mAd041_2 mAd042_1 mAd042_2 mAd043_1 mAd043_2 mAd044_1 mAd044_2 mAd045_1 mAd045_2 mAd046_1 mAd046_2 mAd047_1 mAd047_2 mAd050_1 mAd050_2 mAd051_1 mAd051_2 mAd052_1 mAd052_2 mAd053_1 mAd053_2 mAd054_1 mAd054_2 mAd055_1 mAd055_2 mAd056_1 mAd056_2 mAd057_1 mAd057_2 mAd060_1 mAd060_2 mAd066_1 mAd066_2 mAd067_1 mAd067_2 mAd100_1 mAd100_2 mAd101_1 
+mAd101_2 mAd102_1 mAd102_2 mAd110_1 mAd110_2 mAd111_1 mAd111_2 mAd112_1 mAd112_2 mAd113_1 mAd113_2 mAd114_1 mAd114_2 mAd115_1 mAd115_2 mAd116_1 mAd116_2 mAd117_1 mAd117_2 mAd120_1 mAd120_2 mAd121_1 mAd121_2 mAd122_1 mAd122_2 mAd123_1 mAd123_2 mAd124_1 mAd124_2 mAd125_1 mAd125_2 mAd126_1 mAd126_2 mAd127_1 mAd127_2 mAd130_1 mAd130_2 mAd131_1 mAd131_2 mAd132_1 mAd132_2 mAd133_1 mAd133_2 mAd134_1 mAd134_2 mAd135_1 mAd135_2 mAd136_1 mAd136_2 mAd137_1 mAd137_2 mAd140_1 mAd140_2 mAd141_1 mAd141_2 mAd142_1 
+mAd142_2 mAd143_1 mAd143_2 mAd144_1 mAd144_2 mAd145_1 mAd145_2 mAd146_1 mAd146_2 mAd147_1 mAd147_2 mAd150_1 mAd150_2 mAd151_1 mAd151_2 mAd152_1 mAd152_2 mAd153_1 mAd153_2 mAd154_1 mAd154_2 mAd155_1 mAd155_2 mAd156_1 mAd156_2 mAd157_1 mAd157_2 mAd160_1 mAd160_2 mAd161_1 mAd161_2 mAd162_1 mAd162_2 mAd163_1 mAd163_2 mAd164_1 mAd164_2 mAd165_1 mAd165_2 mAd166_1 mAd166_2 mAd167_1 mAd167_2 mAd170_1 mAd170_2 mAd171_1 mAd171_2 mAd172_1 mAd172_2 mAd173_1 mAd173_2 mAd175_1 mAd175_2 mAd176_1 mAd176_2 mAd177_1 
+mAd177_2 mAd200_1 mAd200_2 mAd201_1 mAd201_2 mAd202_1 mAd202_2 mAd204_1 mAd204_2 mAd205_1 mAd205_2 mAd206_1 mAd206_2 mAd207_1 mAd207_2 mAd210_1 mAd210_2 mAd211_1 mAd211_2 mAd212_1 mAd212_2 mAd213_1 mAd213_2 mAd214_1 mAd214_2 mAd215_1 mAd215_2 mAd216_1 mAd216_2 mAd217_1 mAd217_2 mAd220_1 mAd220_2 mAd221_1 mAd221_2 mAd222_1 mAd222_2 mAd223_1 mAd223_2 mAd224_1 mAd224_2 mAd225_1 mAd225_2 mAd226_1 mAd226_2 mAd227_1 mAd227_2 mAd230_1 mAd230_2 mAd231_1 mAd231_2 mAd232_1 mAd232_2 mAd233_1 mAd233_2 mAd234_1 
+mAd234_2 mAd235_1 mAd235_2 mAd236_1 mAd236_2 mAd237_1 mAd237_2 mAd240_1 mAd240_2 mAd241_1 mAd241_2 mAd242_1 mAd242_2 mAd243_1 mAd243_2 mAd244_1 mAd244_2 mAd245_1 mAd245_2 mAd246_1 mAd246_2 mAd247_1 mAd247_2 mAd250_1 mAd250_2 mAd251_1 mAd251_2 mAd252_1 mAd252_2 mAd253_1 mAd253_2 mAd254_1 mAd254_2 mAd255_1 mAd255_2 mAd256_1 mAd256_2 mAd257_1 mAd257_2 mAd260_1 mAd260_2 mAd261_1 mAd261_2 mAd262_1 mAd262_2 mAd263_1 mAd263_2 mAd264_1 mAd264_2 mAd265_1 mAd265_2 mAd266_1 mAd266_2 mAd267_1 mAd267_2 mAd275_1 
+mAd275_2 mAd276_1 mAd276_2 mAd277_1 mAd277_2 mAd300_1 mAd300_2 mAd310_1 mAd310_2 mAd311_1 mAd311_2 mAd317_1 mAd317_2 mAd320_1 mAd320_2 mAd321_1 mAd321_2 mAd322_1 mAd322_2 mAd323_1 mAd323_2 mAd324_1 mAd324_2 mAd325_1 mAd325_2 mAd326_1 mAd326_2 mAd327_1 mAd327_2 mAd330_1 mAd330_2 mAd331_1 mAd331_2 mAd332_1 mAd332_2 mAd333_1 mAd333_2 mAd334_1 mAd334_2 mAd335_1 mAd335_2 mAd336_1 mAd336_2 mAd337_1 mAd337_2 mAd340_1 mAd340_2 mAd341_1 mAd341_2 mAd342_1 mAd342_2 mAd343_1 mAd343_2 mAd344_1 mAd344_2 mAd345_1 
+mAd345_2 mAd346_1 mAd346_2 mAd347_1 mAd347_2 mAd350_1 mAd350_2 mAd351_1 mAd351_2 mAd352_1 mAd352_2 mAd353_1 mAd353_2 mAd354_1 mAd354_2 mAd355_1 mAd355_2 mAd356_1 mAd356_2 mAd357_1 mAd357_2 mAd360_1 mAd360_2 mAd361_1 mAd361_2 mAd362_1 mAd362_2 mAd363_1 mAd363_2 mAd364_1 mAd364_2 mAd365_1 mAd365_2 mAd366_1 mAd366_2 mAd367_1 mAd367_2 mAd371_1 mAd371_2 mAd372_1 mAd372_2 mAd373_1 mAd373_2 mAd374_1 mAd374_2 mAd375_1 mAd375_2 mAd376_1 mAd376_2 mAd377_1 mAd377_2 mAd400_1 mAd400_2 mAd401_1 mAd401_2 mAd402_1 
+mAd402_2 mAd403_1 mAd403_2 mAd404_1 mAd404_2 mAd405_1 mAd405_2 mAd406_1 mAd406_2 mAd407_1 mAd407_2 mAd410_1 mAd410_2 mAd411_1 mAd411_2 mAd412_1 mAd412_2 mAd413_1 mAd413_2 mAd414_1 mAd414_2 mAd415_1 mAd415_2 mAd416_1 mAd416_2 mAd417_1 mAd417_2 mAd420_1 mAd420_2 mAd421_1 mAd421_2 mAd422_1 mAd422_2 mAd423_1 mAd423_2 mAd424_1 mAd424_2 mAd425_1 mAd425_2 mAd426_1 mAd426_2 mAd427_1 mAd427_2 mAd430_1 mAd430_2 mAd431_1 mAd431_2 mAd432_1 mAd432_2 mAd433_1 mAd433_2 mAd434_1 mAd434_2 mAd435_1 mAd435_2 mAd436_1 
+mAd436_2 mAd437_1 mAd437_2 mAd440_1 mAd440_2 mAd441_1 mAd441_2 mAd442_1 mAd442_2 mAd443_1 mAd443_2 mAd444_1 mAd444_2 mAd445_1 mAd445_2 mAd446_1 mAd446_2 mAd447_1 mAd447_2 mAd450_1 mAd450_2 mAd451_1 mAd451_2 mAd452_1 mAd452_2 mAd453_1 mAd453_2 mAd454_1 mAd454_2 mAd455_1 mAd455_2 mAd456_1 mAd456_2 mAd457_1 mAd457_2 mAd460_1 mAd460_2 mAd466_1 mAd466_2 mAd467_1 mAd467_2 mAd500_1 mAd500_2 mAd501_1 mAd501_2 mAd502_1 mAd502_2 mAd508_1 mAd508_2 mAd509_1 mAd509_2 mAd512_1 mAd512_2 mAd513_1 mAd513_2 mAd514_1 
+mAd514_2 mAd515_1 mAd515_2 mAd516_1 mAd516_2 mAd517_1 mAd517_2 mAd520_1 mAd520_2 mAd521_1 mAd521_2 mAd522_1 mAd522_2 mAd523_1 mAd523_2 mAd524_1 mAd524_2 mAd525_1 mAd525_2 mAd526_1 mAd526_2 mAd527_1 mAd527_2 mAd530_1 mAd530_2 mAd531_1 mAd531_2 mAd532_1 mAd532_2 mAd533_1 mAd533_2 mAd534_1 mAd534_2 mAd535_1 mAd535_2 mAd536_1 mAd536_2 mAd537_1 mAd537_2 mAd540_1 mAd540_2 mAd541_1 mAd541_2 mAd542_1 mAd542_2 mAd543_1 mAd543_2 mAd544_1 mAd544_2 mAd545_1 mAd545_2 mAd546_1 mAd546_2 mAd547_1 mAd547_2 mAd550_1 
+mAd550_2 mAd551_1 mAd551_2 mAd552_1 mAd552_2 mAd553_1 mAd553_2 mAd554_1 mAd554_2 mAd555_1 mAd555_2 mAd556_1 mAd556_2 mAd557_1 mAd557_2 mAd560_1 mAd560_2 mAd561_1 mAd561_2 mAd562_1 mAd562_2 mAd563_1 mAd563_2 mAd564_1 mAd564_2 mAd565_1 mAd565_2 mAd566_1 mAd566_2 mAd567_1 mAd567_2 mAd570_1 mAd570_2 mAd571_1 mAd571_2 mAd572_1 mAd572_2 mAd573_1 mAd573_2 mAd575_1 mAd575_2 mAd576_1 mAd576_2 mAd577_1 mAd577_2 mAd600_1 mAd600_2 mAd601_1 mAd601_2 mAd602_1 mAd602_2 mAd604_1 mAd604_2 mAd605_1 mAd605_2 mAd606_1 
+mAd606_2 mAd607_1 mAd607_2 mAd610_1 mAd610_2 mAd611_1 mAd611_2 mAd612_1 mAd612_2 mAd613_1 mAd613_2 mAd614_1 mAd614_2 mAd615_1 mAd615_2 mAd616_1 mAd616_2 mAd617_1 mAd617_2 mAd620_1 mAd620_2 mAd621_1 mAd621_2 mAd622_1 mAd622_2 mAd623_1 mAd623_2 mAd624_1 mAd624_2 mAd625_1 mAd625_2 mAd626_1 mAd626_2 mAd627_1 mAd627_2 mAd630_1 mAd630_2 mAd631_1 mAd631_2 mAd632_1 mAd632_2 mAd633_1 mAd633_2 mAd634_1 mAd634_2 mAd635_1 mAd635_2 mAd636_1 mAd636_2 mAd637_1 mAd637_2 mAd640_1 mAd640_2 mAd641_1 mAd641_2 mAd642_1 
+mAd642_2 mAd643_1 mAd643_2 mAd644_1 mAd644_2 mAd645_1 mAd645_2 mAd646_1 mAd646_2 mAd647_1 mAd647_2 mAd650_1 mAd650_2 mAd651_1 mAd651_2 mAd652_1 mAd652_2 mAd653_1 mAd653_2 mAd654_1 mAd654_2 mAd655_1 mAd655_2 mAd656_1 mAd656_2 mAd657_1 mAd657_2 mAd660_1 mAd660_2 mAd661_1 mAd661_2 mAd662_1 mAd662_2 mAd663_1 mAd663_2 mAd664_1 mAd664_2 mAd665_1 mAd665_2 mAd666_1 mAd666_2 mAd667_1 mAd667_2 mAd675_1 mAd675_2 mAd676_1 mAd676_2 mAd677_1 mAd677_2 mAd700_1 mAd700_2 mAd710_1 mAd710_2 mAd711_1 mAd711_2 mAd717_1 
+mAd717_2 mAd720_1 mAd720_2 mAd721_1 mAd721_2 mAd722_1 mAd722_2 mAd723_1 mAd723_2 mAd724_1 mAd724_2 mAd725_1 mAd725_2 mAd726_1 mAd726_2 mAd727_1 mAd727_2 mAd730_1 mAd730_2 mAd731_1 mAd731_2 mAd732_1 mAd732_2 mAd733_1 mAd733_2 mAd734_1 mAd734_2 mAd735_1 mAd735_2 mAd736_1 mAd736_2 mAd737_1 mAd737_2 mAd740_1 mAd740_2 mAd741_1 mAd741_2 mAd742_1 mAd742_2 mAd743_1 mAd743_2 mAd744_1 mAd744_2 mAd745_1 mAd745_2 mAd746_1 mAd746_2 mAd747_1 mAd747_2 mAd750_1 mAd750_2 mAd751_1 mAd751_2 mAd752_1 mAd752_2 mAd753_1 
+mAd753_2 mAd754_1 mAd754_2 mAd755_1 mAd755_2 mAd756_1 mAd756_2 mAd757_1 mAd757_2 mAd760_1 mAd760_2 mAd761_1 mAd761_2 mAd762_1 mAd762_2 mAd763_1 mAd763_2 mAd764_1 mAd764_2 mAd765_1 mAd765_2 mAd766_1 mAd766_2 mAd767_1 mAd767_2 mAd771_1 mAd771_2 mAd772_1 mAd772_2 mAd773_1 mAd773_2 mAd774_1 mAd774_2 mAd775_1 mAd775_2 mAd776_1 mAd776_2 mAd777_1 mAd777_2 X0 X1 X10 X11 X12 X13 X2 X3 X4 X5 X6 X7 X8 X9 Y1 Y10 Y11 Y12 Y2 Y3 Y4 Y5 Y6 Y7 Y8 Y9 Z1 Z10 Z11 Z12 Z2 Z3 Z4 Z5 Z6 Z7 Z8 Z9
** GLOBAL gnd
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
Xkey@3 mAd067_1 mAd067_2 K0 X0 basic__key adr=67
Xkey@4 mAd056_1 mAd056_2 X1 Y1 basic__key adr=56
Xkey@5 mAd054_1 mAd054_2 Y1 a2 basic__key adr=54
Xkey@6 mAd046_1 mAd046_2 X1 a1 basic__key adr=46
Xkey@8 mAd044_1 mAd044_2 a1 a2 basic__key adr=44
Xkey@9 mAd055_1 mAd055_2 X1 a2 basic__key adr=55
Xkey@10 mAd045_1 mAd045_2 Y1 a1 basic__key adr=45
Xkey@11 mAd066_1 mAd066_2 Y1 X0 basic__key adr=66
Xkey@12 mAd057_1 mAd057_2 K0 X1 basic__key adr=57
Xkey@13 mAd323_1 mAd323_2 a6 Y12 basic__key adr=323
Xkey@14 mAd321_1 mAd321_2 Y12 Z1 basic__key adr=321
Xkey@15 mAd333_1 mAd333_2 a6 a7 basic__key adr=333
Xkey@16 mAd331_1 mAd331_2 a7 Z1 basic__key adr=331
Xkey@17 mAd322_1 mAd322_2 a6 Z1 basic__key adr=322
Xkey@18 mAd332_1 mAd332_2 Y12 a7 basic__key adr=332
Xkey@19 mAd121_1 mAd121_2 a2 Y6 basic__key adr=121
Xkey@20 mAd160_1 mAd160_2 Y6 a4 basic__key adr=160
Xkey@21 mAd111_1 mAd111_2 a2 a3 basic__key adr=111
Xkey@22 mAd150_1 mAd150_2 a3 a4 basic__key adr=150
Xkey@23 mAd100_1 mAd100_2 a2 a4 basic__key adr=100
Xkey@24 mAd171_1 mAd171_2 Y6 a3 basic__key adr=171
Xkey@25 mAd217_1 mAd217_2 a4 Y7 basic__key adr=217
Xkey@26 mAd256_1 mAd256_2 Y7 a6 basic__key adr=256
Xkey@27 mAd227_1 mAd227_2 a4 a5 basic__key adr=227
Xkey@28 mAd266_1 mAd266_2 a5 a6 basic__key adr=266
Xkey@29 mAd277_1 mAd277_2 a4 a6 basic__key adr=277
Xkey@30 mAd206_1 mAd206_2 Y7 a5 basic__key adr=206
Xkey@31 mAd035_1 mAd035_2 X2 Y2 basic__key adr=35
Xkey@32 mAd033_1 mAd033_2 Y2 b2 basic__key adr=33
Xkey@33 mAd025_1 mAd025_2 X2 b1 basic__key adr=25
Xkey@34 mAd023_1 mAd023_2 b1 b2 basic__key adr=23
Xkey@35 mAd034_1 mAd034_2 X2 b2 basic__key adr=34
Xkey@36 mAd024_1 mAd024_2 Y2 b1 basic__key adr=24
Xkey@37 mAd014_1 mAd014_2 X3 Y3 basic__key adr=14
Xkey@38 mAd012_1 mAd012_2 Y3 c2 basic__key adr=12
Xkey@39 mAd004_1 mAd004_2 X3 c1 basic__key adr=4
Xkey@40 mAd002_1 mAd002_2 c1 c2 basic__key adr=2
Xkey@41 mAd013_1 mAd013_2 X3 c2 basic__key adr=13
Xkey@42 mAd003_1 mAd003_2 Y3 c1 basic__key adr=3
Xkey@43 mAd126_1 mAd126_2 d2 c3 basic__key adr=126
Xkey@44 mAd124_1 mAd124_2 c3 d4 basic__key adr=124
Xkey@45 mAd116_1 mAd116_2 d2 d3 basic__key adr=116
Xkey@46 mAd114_1 mAd114_2 d3 d4 basic__key adr=114
Xkey@47 mAd125_1 mAd125_2 d2 d4 basic__key adr=125
Xkey@48 mAd115_1 mAd115_2 c3 d3 basic__key adr=115
Xkey@49 mAd145_1 mAd145_2 e2 b3 basic__key adr=145
Xkey@50 mAd143_1 mAd143_2 b3 e4 basic__key adr=143
Xkey@51 mAd135_1 mAd135_2 e2 e3 basic__key adr=135
Xkey@52 mAd133_1 mAd133_2 e3 e4 basic__key adr=133
Xkey@53 mAd144_1 mAd144_2 e2 e4 basic__key adr=144
Xkey@54 mAd134_1 mAd134_2 b3 e3 basic__key adr=134
Xkey@55 mAd164_1 mAd164_2 f2 a3 basic__key adr=164
Xkey@56 mAd142_1 mAd142_2 a3 f4 basic__key adr=142
Xkey@57 mAd154_1 mAd154_2 f2 f3 basic__key adr=154
Xkey@58 mAd132_1 mAd132_2 f3 f4 basic__key adr=132
Xkey@59 mAd163_1 mAd163_2 f2 f4 basic__key adr=163
Xkey@60 mAd153_1 mAd153_2 a3 f3 basic__key adr=153
Xkey@61 mAd645_1 mAd645_2 g4 f5 basic__key adr=645
Xkey@62 mAd623_1 mAd623_2 f5 g6 basic__key adr=623
Xkey@63 mAd635_1 mAd635_2 g4 g5 basic__key adr=635
Xkey@64 mAd613_1 mAd613_2 g5 g6 basic__key adr=613
Xkey@65 mAd614_1 mAd614_2 g4 g6 basic__key adr=614
Xkey@66 mAd624_1 mAd624_2 f5 g5 basic__key adr=624
Xkey@67 mAd644_1 mAd644_2 h4 e5 basic__key adr=644
Xkey@68 mAd642_1 mAd642_2 e5 h6 basic__key adr=642
Xkey@69 mAd634_1 mAd634_2 h4 h5 basic__key adr=634
Xkey@70 mAd632_1 mAd632_2 h5 h6 basic__key adr=632
Xkey@71 mAd633_1 mAd633_2 h4 h6 basic__key adr=633
Xkey@72 mAd643_1 mAd643_2 e5 h5 basic__key adr=643
Xkey@73 mAd663_1 mAd663_2 i4 d5 basic__key adr=663
Xkey@74 mAd661_1 mAd661_2 d5 i6 basic__key adr=661
Xkey@75 mAd653_1 mAd653_2 i4 i5 basic__key adr=653
Xkey@76 mAd651_1 mAd651_2 i5 i6 basic__key adr=651
Xkey@77 mAd652_1 mAd652_2 i4 i6 basic__key adr=652
Xkey@78 mAd662_1 mAd662_2 d5 i5 basic__key adr=662
Xkey@79 mAd775_1 mAd775_2 j3 i7 basic__key adr=775
Xkey@80 mAd773_1 mAd773_2 i7 Z10 basic__key adr=773
Xkey@81 mAd765_1 mAd765_2 j3 K10 basic__key adr=765
Xkey@82 mAd763_1 mAd763_2 K10 Z10 basic__key adr=763
Xkey@83 mAd764_1 mAd764_2 j3 Z10 basic__key adr=764
Xkey@84 mAd774_1 mAd774_2 i7 K10 basic__key adr=774
Xkey@85 mAd754_1 mAd754_2 k3 h7 basic__key adr=754
Xkey@86 mAd752_1 mAd752_2 h7 Z11 basic__key adr=752
Xkey@87 mAd744_1 mAd744_2 k3 K11 basic__key adr=744
Xkey@88 mAd742_1 mAd742_2 K11 Z11 basic__key adr=742
Xkey@89 mAd743_1 mAd743_2 k3 Z11 basic__key adr=743
Xkey@90 mAd753_1 mAd753_2 h7 K11 basic__key adr=753
Xkey@91 mAd733_1 mAd733_2 l3 g7 basic__key adr=733
Xkey@92 mAd731_1 mAd731_2 g7 Z12 basic__key adr=731
Xkey@93 mAd723_1 mAd723_2 l3 K12 basic__key adr=723
Xkey@94 mAd721_1 mAd721_2 K12 Z12 basic__key adr=721
Xkey@95 mAd722_1 mAd722_2 l3 Z12 basic__key adr=722
Xkey@96 mAd732_1 mAd732_2 g7 K12 basic__key adr=732
Xkey@97 mAd037_1 mAd037_2 K0 X2 basic__key adr=37
Xkey@98 mAd017_1 mAd017_2 K0 X3 basic__key adr=17
Xkey@99 mAd007_1 mAd007_2 K0 X4 basic__key adr=7
Xkey@100 mAd027_1 mAd027_2 K0 X5 basic__key adr=27
Xkey@101 mAd047_1 mAd047_2 K0 X6 basic__key adr=47
Xkey@102 mAd447_1 mAd447_2 K0 X7 basic__key adr=447
Xkey@103 mAd427_1 mAd427_2 K0 X8 basic__key adr=427
Xkey@104 mAd407_1 mAd407_2 K0 X9 basic__key adr=407
Xkey@105 mAd417_1 mAd417_2 K0 X10 basic__key adr=417
Xkey@106 mAd437_1 mAd437_2 K0 X11 basic__key adr=437
Xkey@107 mAd457_1 mAd457_2 K0 X12 basic__key adr=457
Xkey@108 mAd467_1 mAd467_2 K0 X13 basic__key adr=467
Xkey@109 mAd446_1 mAd446_2 X12 g1 basic__key adr=446
Xkey@110 mAd444_1 mAd444_2 g1 l1 basic__key adr=444
Xkey@111 mAd456_1 mAd456_2 X12 K1 basic__key adr=456
Xkey@112 mAd454_1 mAd454_2 K1 l1 basic__key adr=454
Xkey@113 mAd455_1 mAd455_2 X12 l1 basic__key adr=455
Xkey@114 mAd445_1 mAd445_2 g1 K1 basic__key adr=445
Xkey@115 mAd425_1 mAd425_2 X11 h1 basic__key adr=425
Xkey@116 mAd423_1 mAd423_2 h1 k1 basic__key adr=423
Xkey@117 mAd435_1 mAd435_2 X11 K2 basic__key adr=435
Xkey@118 mAd433_1 mAd433_2 K2 k1 basic__key adr=433
Xkey@119 mAd434_1 mAd434_2 X11 k1 basic__key adr=434
Xkey@120 mAd424_1 mAd424_2 h1 K2 basic__key adr=424
Xkey@121 mAd404_1 mAd404_2 X10 i1 basic__key adr=404
Xkey@122 mAd402_1 mAd402_2 i1 j1 basic__key adr=402
Xkey@123 mAd414_1 mAd414_2 X10 K3 basic__key adr=414
Xkey@124 mAd412_1 mAd412_2 K3 j1 basic__key adr=412
Xkey@125 mAd413_1 mAd413_2 X10 j1 basic__key adr=413
Xkey@126 mAd403_1 mAd403_2 i1 K3 basic__key adr=403
Xkey@127 mAd516_1 mAd516_2 i2 d3 basic__key adr=516
Xkey@128 mAd514_1 mAd514_2 d3 i4 basic__key adr=514
Xkey@129 mAd526_1 mAd526_2 i2 i3 basic__key adr=526
Xkey@130 mAd524_1 mAd524_2 i3 i4 basic__key adr=524
Xkey@131 mAd525_1 mAd525_2 i2 i4 basic__key adr=525
Xkey@132 mAd515_1 mAd515_2 d3 i3 basic__key adr=515
Xkey@133 mAd535_1 mAd535_2 h2 e3 basic__key adr=535
Xkey@134 mAd533_1 mAd533_2 e3 h4 basic__key adr=533
Xkey@135 mAd545_1 mAd545_2 h2 h3 basic__key adr=545
Xkey@136 mAd543_1 mAd543_2 h3 h4 basic__key adr=543
Xkey@137 mAd544_1 mAd544_2 h2 h4 basic__key adr=544
Xkey@138 mAd534_1 mAd534_2 e3 h3 basic__key adr=534
Xkey@139 mAd554_1 mAd554_2 g2 f3 basic__key adr=554
Xkey@140 mAd532_1 mAd532_2 f3 g4 basic__key adr=532
Xkey@141 mAd564_1 mAd564_2 g2 g3 basic__key adr=564
Xkey@142 mAd542_1 mAd542_2 g3 g4 basic__key adr=542
Xkey@143 mAd563_1 mAd563_2 g2 g4 basic__key adr=563
Xkey@144 mAd553_1 mAd553_2 f3 g3 basic__key adr=553
Xkey@145 mAd235_1 mAd235_2 f4 a5 basic__key adr=235
Xkey@146 mAd213_1 mAd213_2 a5 f6 basic__key adr=213
Xkey@147 mAd245_1 mAd245_2 f4 f5 basic__key adr=245
Xkey@148 mAd223_1 mAd223_2 f5 f6 basic__key adr=223
Xkey@149 mAd214_1 mAd214_2 f4 f6 basic__key adr=214
Xkey@150 mAd224_1 mAd224_2 a5 f5 basic__key adr=224
Xkey@151 mAd234_1 mAd234_2 e4 b5 basic__key adr=234
Xkey@152 mAd232_1 mAd232_2 b5 e6 basic__key adr=232
Xkey@153 mAd244_1 mAd244_2 e4 e5 basic__key adr=244
Xkey@154 mAd242_1 mAd242_2 e5 e6 basic__key adr=242
Xkey@155 mAd233_1 mAd233_2 e4 e6 basic__key adr=233
Xkey@156 mAd243_1 mAd243_2 b5 e5 basic__key adr=243
Xkey@157 mAd253_1 mAd253_2 d4 c5 basic__key adr=253
Xkey@158 mAd251_1 mAd251_2 c5 d6 basic__key adr=251
Xkey@159 mAd263_1 mAd263_2 d4 d5 basic__key adr=263
Xkey@160 mAd261_1 mAd261_2 d5 d6 basic__key adr=261
Xkey@161 mAd252_1 mAd252_2 d4 d6 basic__key adr=252
Xkey@162 mAd262_1 mAd262_2 c5 d5 basic__key adr=262
Xkey@163 mAd365_1 mAd365_2 c6 Y10 basic__key adr=365
Xkey@164 mAd363_1 mAd363_2 Y10 Z3 basic__key adr=363
Xkey@165 mAd375_1 mAd375_2 c6 c7 basic__key adr=375
Xkey@166 mAd373_1 mAd373_2 c7 Z3 basic__key adr=373
Xkey@167 mAd364_1 mAd364_2 c6 Z3 basic__key adr=364
Xkey@168 mAd374_1 mAd374_2 Y10 c7 basic__key adr=374
Xkey@169 mAd344_1 mAd344_2 b6 Y11 basic__key adr=344
Xkey@170 mAd342_1 mAd342_2 Y11 Z2 basic__key adr=342
Xkey@171 mAd354_1 mAd354_2 b6 b7 basic__key adr=354
Xkey@172 mAd352_1 mAd352_2 b7 Z2 basic__key adr=352
Xkey@173 mAd343_1 mAd343_2 b6 Z2 basic__key adr=343
Xkey@174 mAd353_1 mAd353_2 Y11 b7 basic__key adr=353
Xkey@175 mAd122_1 mAd122_2 b2 Y5 basic__key adr=122
Xkey@176 mAd161_1 mAd161_2 Y5 b4 basic__key adr=161
Xkey@177 mAd112_1 mAd112_2 b2 b3 basic__key adr=112
Xkey@178 mAd151_1 mAd151_2 b3 b4 basic__key adr=151
Xkey@179 mAd101_1 mAd101_2 b2 b4 basic__key adr=101
Xkey@180 mAd172_1 mAd172_2 Y5 b3 basic__key adr=172
Xkey@181 mAd123_1 mAd123_2 c2 Y4 basic__key adr=123
Xkey@182 mAd162_1 mAd162_2 Y4 c4 basic__key adr=162
Xkey@183 mAd113_1 mAd113_2 c2 c3 basic__key adr=113
Xkey@184 mAd152_1 mAd152_2 c3 c4 basic__key adr=152
Xkey@185 mAd102_1 mAd102_2 c2 c4 basic__key adr=102
Xkey@186 mAd173_1 mAd173_2 Y4 c3 basic__key adr=173
Xkey@187 mAd011_1 mAd011_2 X4 c1 basic__key adr=11
Xkey@188 mAd127_1 mAd127_2 c1 d2 basic__key adr=127
Xkey@189 mAd001_1 mAd001_2 X4 d1 basic__key adr=1
Xkey@190 mAd117_1 mAd117_2 d1 d2 basic__key adr=117
Xkey@191 mAd010_1 mAd010_2 X4 d2 basic__key adr=10
Xkey@192 mAd000_1 mAd000_2 c1 d1 basic__key adr=0
Xkey@193 mAd032_1 mAd032_2 X5 b1 basic__key adr=32
Xkey@194 mAd030_1 mAd030_2 b1 e2 basic__key adr=30
Xkey@195 mAd022_1 mAd022_2 X5 e1 basic__key adr=22
Xkey@196 mAd020_1 mAd020_2 e1 e2 basic__key adr=20
Xkey@197 mAd031_1 mAd031_2 X5 e2 basic__key adr=31
Xkey@198 mAd021_1 mAd021_2 b1 e1 basic__key adr=21
Xkey@199 mAd053_1 mAd053_2 X6 a1 basic__key adr=53
Xkey@200 mAd051_1 mAd051_2 a1 f2 basic__key adr=51
Xkey@201 mAd043_1 mAd043_2 X6 f1 basic__key adr=43
Xkey@202 mAd041_1 mAd041_2 f1 f2 basic__key adr=41
Xkey@203 mAd052_1 mAd052_2 X6 f2 basic__key adr=52
Xkey@204 mAd042_1 mAd042_2 a1 f1 basic__key adr=42
Xkey@205 mAd443_1 mAd443_2 X7 f1 basic__key adr=443
Xkey@206 mAd441_1 mAd441_2 f1 g2 basic__key adr=441
Xkey@207 mAd453_1 mAd453_2 X7 g1 basic__key adr=453
Xkey@208 mAd451_1 mAd451_2 g1 g2 basic__key adr=451
Xkey@209 mAd452_1 mAd452_2 X7 g2 basic__key adr=452
Xkey@210 mAd442_1 mAd442_2 f1 g1 basic__key adr=442
Xkey@211 mAd422_1 mAd422_2 X8 e1 basic__key adr=422
Xkey@212 mAd420_1 mAd420_2 e1 h2 basic__key adr=420
Xkey@213 mAd432_1 mAd432_2 X8 h1 basic__key adr=432
Xkey@214 mAd430_1 mAd430_2 h1 h2 basic__key adr=430
Xkey@215 mAd431_1 mAd431_2 X8 h2 basic__key adr=431
Xkey@216 mAd421_1 mAd421_2 e1 h1 basic__key adr=421
Xkey@217 mAd401_1 mAd401_2 X9 d1 basic__key adr=401
Xkey@218 mAd517_1 mAd517_2 d1 i2 basic__key adr=517
Xkey@219 mAd411_1 mAd411_2 X9 i1 basic__key adr=411
Xkey@220 mAd527_1 mAd527_2 i1 i2 basic__key adr=527
Xkey@221 mAd410_1 mAd410_2 X9 i2 basic__key adr=410
Xkey@222 mAd400_1 mAd400_2 d1 i1 basic__key adr=400
Xkey@223 mAd513_1 mAd513_2 j1 i3 basic__key adr=513
Xkey@224 mAd552_1 mAd552_2 i3 j2 basic__key adr=552
Xkey@225 mAd523_1 mAd523_2 j1 K4 basic__key adr=523
Xkey@226 mAd562_1 mAd562_2 K4 j2 basic__key adr=562
Xkey@227 mAd502_1 mAd502_2 j1 j2 basic__key adr=502
Xkey@228 mAd573_1 mAd573_2 i3 K4 basic__key adr=573
Xkey@229 mAd512_1 mAd512_2 k1 h3 basic__key adr=512
Xkey@230 mAd551_1 mAd551_2 h3 k2 basic__key adr=551
Xkey@231 mAd522_1 mAd522_2 k1 K5 basic__key adr=522
Xkey@232 mAd561_1 mAd561_2 K5 k2 basic__key adr=561
Xkey@233 mAd501_1 mAd501_2 k1 k2 basic__key adr=501
Xkey@234 mAd572_1 mAd572_2 h3 K5 basic__key adr=572
Xkey@235 mAd509_1 mAd509_2 l1 g3 basic__key adr=509
Xkey@236 mAd550_1 mAd550_2 g3 l2 basic__key adr=550
Xkey@237 mAd521_1 mAd521_2 l1 K6 basic__key adr=521
Xkey@238 mAd560_1 mAd560_2 K6 l2 basic__key adr=560
Xkey@239 mAd500_1 mAd500_2 l1 l2 basic__key adr=500
Xkey@240 mAd571_1 mAd571_2 g3 K6 basic__key adr=571
Xkey@241 mAd627_1 mAd627_2 l2 g5 basic__key adr=627
Xkey@242 mAd666_1 mAd666_2 g5 l3 basic__key adr=666
Xkey@243 mAd617_1 mAd617_2 l2 K7 basic__key adr=617
Xkey@244 mAd656_1 mAd656_2 K7 l3 basic__key adr=656
Xkey@245 mAd677_1 mAd677_2 l2 l3 basic__key adr=677
Xkey@246 mAd606_1 mAd606_2 g5 K7 basic__key adr=606
Xkey@247 mAd626_1 mAd626_2 k2 h5 basic__key adr=626
Xkey@248 mAd665_1 mAd665_2 h5 k3 basic__key adr=665
Xkey@249 mAd616_1 mAd616_2 k2 K8 basic__key adr=616
Xkey@250 mAd655_1 mAd655_2 K8 k3 basic__key adr=655
Xkey@251 mAd676_1 mAd676_2 k2 k3 basic__key adr=676
Xkey@252 mAd605_1 mAd605_2 h5 K8 basic__key adr=605
Xkey@253 mAd625_1 mAd625_2 j2 i5 basic__key adr=625
Xkey@254 mAd664_1 mAd664_2 i5 j3 basic__key adr=664
Xkey@255 mAd615_1 mAd615_2 j2 K9 basic__key adr=615
Xkey@256 mAd654_1 mAd654_2 K9 j3 basic__key adr=654
Xkey@257 mAd675_1 mAd675_2 j2 j3 basic__key adr=675
Xkey@258 mAd604_1 mAd604_2 i5 K9 basic__key adr=604
Xkey@259 mAd660_1 mAd660_2 i6 d7 basic__key adr=660
Xkey@260 mAd776_1 mAd776_2 d7 Z9 basic__key adr=776
Xkey@261 mAd650_1 mAd650_2 i6 i7 basic__key adr=650
Xkey@262 mAd766_1 mAd766_2 i7 Z9 basic__key adr=766
Xkey@263 mAd767_1 mAd767_2 i6 Z9 basic__key adr=767
Xkey@264 mAd777_1 mAd777_2 d7 i7 basic__key adr=777
Xkey@265 mAd757_1 mAd757_2 h6 e7 basic__key adr=757
Xkey@266 mAd755_1 mAd755_2 e7 Z8 basic__key adr=755
Xkey@267 mAd747_1 mAd747_2 h6 h7 basic__key adr=747
Xkey@268 mAd745_1 mAd745_2 h7 Z8 basic__key adr=745
Xkey@269 mAd746_1 mAd746_2 h6 Z8 basic__key adr=746
Xkey@270 mAd756_1 mAd756_2 e7 h7 basic__key adr=756
Xkey@271 mAd736_1 mAd736_2 g6 f7 basic__key adr=736
Xkey@272 mAd734_1 mAd734_2 f7 Z7 basic__key adr=734
Xkey@273 mAd726_1 mAd726_2 g6 g7 basic__key adr=726
Xkey@274 mAd724_1 mAd724_2 g7 Z7 basic__key adr=724
Xkey@275 mAd725_1 mAd725_2 g6 Z7 basic__key adr=725
Xkey@276 mAd735_1 mAd735_2 f7 g7 basic__key adr=735
Xkey@277 mAd326_1 mAd326_2 f6 a7 basic__key adr=326
Xkey@278 mAd324_1 mAd324_2 a7 Z6 basic__key adr=324
Xkey@279 mAd336_1 mAd336_2 f6 f7 basic__key adr=336
Xkey@280 mAd334_1 mAd334_2 f7 Z6 basic__key adr=334
Xkey@281 mAd325_1 mAd325_2 f6 Z6 basic__key adr=325
Xkey@282 mAd335_1 mAd335_2 a7 f7 basic__key adr=335
Xkey@283 mAd347_1 mAd347_2 e6 b7 basic__key adr=347
Xkey@284 mAd345_1 mAd345_2 b7 Z5 basic__key adr=345
Xkey@285 mAd357_1 mAd357_2 e6 e7 basic__key adr=357
Xkey@286 mAd355_1 mAd355_2 e7 Z5 basic__key adr=355
Xkey@287 mAd346_1 mAd346_2 e6 Z5 basic__key adr=346
Xkey@288 mAd356_1 mAd356_2 b7 e7 basic__key adr=356
Xkey@289 mAd250_1 mAd250_2 d6 c7 basic__key adr=250
Xkey@290 mAd366_1 mAd366_2 c7 Z4 basic__key adr=366
Xkey@291 mAd260_1 mAd260_2 d6 d7 basic__key adr=260
Xkey@292 mAd376_1 mAd376_2 d7 Z4 basic__key adr=376
Xkey@293 mAd367_1 mAd367_2 d6 Z4 basic__key adr=367
Xkey@294 mAd377_1 mAd377_2 c7 d7 basic__key adr=377
Xkey@295 mAd215_1 mAd215_2 c4 Y9 basic__key adr=215
Xkey@296 mAd254_1 mAd254_2 Y9 c6 basic__key adr=254
Xkey@297 mAd225_1 mAd225_2 c4 c5 basic__key adr=225
Xkey@298 mAd264_1 mAd264_2 c5 c6 basic__key adr=264
Xkey@299 mAd275_1 mAd275_2 c4 c6 basic__key adr=275
Xkey@300 mAd204_1 mAd204_2 Y9 c5 basic__key adr=204
Xkey@301 mAd216_1 mAd216_2 b4 Y8 basic__key adr=216
Xkey@302 mAd255_1 mAd255_2 Y8 b6 basic__key adr=255
Xkey@303 mAd226_1 mAd226_2 b4 b5 basic__key adr=226
Xkey@304 mAd265_1 mAd265_2 b5 b6 basic__key adr=265
Xkey@305 mAd276_1 mAd276_2 b4 b6 basic__key adr=276
Xkey@306 mAd205_1 mAd205_2 Y8 b5 basic__key adr=205
Xkey@307 mAd060_1 mAd060_2 Y2 X0 basic__key adr=60
Xkey@308 mAd177_1 mAd177_2 Y3 X0 basic__key adr=177
Xkey@309 mAd176_1 mAd176_2 Y4 X0 basic__key adr=176
Xkey@310 mAd175_1 mAd175_2 Y5 X0 basic__key adr=175
Xkey@311 mAd170_1 mAd170_2 Y6 X0 basic__key adr=170
Xkey@312 mAd207_1 mAd207_2 Y7 X0 basic__key adr=207
Xkey@313 mAd202_1 mAd202_2 Y8 X0 basic__key adr=202
Xkey@314 mAd201_1 mAd201_2 Y9 X0 basic__key adr=201
Xkey@315 mAd200_1 mAd200_2 Y10 X0 basic__key adr=200
Xkey@316 mAd317_1 mAd317_2 Y11 X0 basic__key adr=317
Xkey@317 mAd311_1 mAd311_2 Y12 X0 basic__key adr=311
Xkey@318 mAd300_1 mAd300_2 K13 X0 basic__key adr=300
Xkey@319 mAd050_1 mAd050_2 Y2 a2 basic__key adr=50
Xkey@320 mAd167_1 mAd167_2 Y3 a2 basic__key adr=167
Xkey@321 mAd166_1 mAd166_2 Y4 a2 basic__key adr=166
Xkey@322 mAd165_1 mAd165_2 Y5 a2 basic__key adr=165
Xkey@323 mAd212_1 mAd212_2 Y8 a6 basic__key adr=212
Xkey@324 mAd211_1 mAd211_2 Y9 a6 basic__key adr=211
Xkey@325 mAd210_1 mAd210_2 Y10 a6 basic__key adr=210
Xkey@326 mAd327_1 mAd327_2 Y11 a6 basic__key adr=327
Xkey@327 mAd310_1 mAd310_2 K13 Z1 basic__key adr=310
Xkey@328 mAd036_1 mAd036_2 a1 X2 basic__key adr=36
Xkey@329 mAd147_1 mAd147_2 Y3 b2 basic__key adr=147
Xkey@330 mAd146_1 mAd146_2 Y4 b2 basic__key adr=146
Xkey@331 mAd140_1 mAd140_2 a3 b4 basic__key adr=140
Xkey@332 mAd237_1 mAd237_2 a5 b4 basic__key adr=237
Xkey@333 mAd231_1 mAd231_2 Y9 b6 basic__key adr=231
Xkey@334 mAd230_1 mAd230_2 Y10 b6 basic__key adr=230
Xkey@335 mAd341_1 mAd341_2 a7 Z2 basic__key adr=341
Xkey@336 mAd330_1 mAd330_2 K13 Z2 basic__key adr=330
Xkey@337 mAd016_1 mAd016_2 a1 X3 basic__key adr=16
Xkey@338 mAd015_1 mAd015_2 b1 X3 basic__key adr=15
Xkey@339 mAd141_1 mAd141_2 b3 c4 basic__key adr=141
Xkey@340 mAd120_1 mAd120_2 a3 c4 basic__key adr=120
Xkey@341 mAd257_1 mAd257_2 a5 c4 basic__key adr=257
Xkey@342 mAd236_1 mAd236_2 b5 c4 basic__key adr=236
Xkey@343 mAd362_1 mAd362_2 b7 Z3 basic__key adr=362
Xkey@344 mAd361_1 mAd361_2 a7 Z3 basic__key adr=361
Xkey@345 mAd350_1 mAd350_2 K13 Z3 basic__key adr=350
Xkey@346 mAd360_1 mAd360_2 K13 Z4 basic__key adr=360
Xkey@347 mAd371_1 mAd371_2 a7 Z4 basic__key adr=371
Xkey@348 mAd372_1 mAd372_2 b7 Z4 basic__key adr=372
Xkey@349 mAd246_1 mAd246_2 b5 d4 basic__key adr=246
Xkey@350 mAd267_1 mAd267_2 a5 d4 basic__key adr=267
Xkey@351 mAd110_1 mAd110_2 a3 d4 basic__key adr=110
Xkey@352 mAd131_1 mAd131_2 b3 d4 basic__key adr=131
Xkey@353 mAd005_1 mAd005_2 b1 X4 basic__key adr=5
Xkey@354 mAd006_1 mAd006_2 a1 X4 basic__key adr=6
Xkey@355 mAd026_1 mAd026_2 a1 X5 basic__key adr=26
Xkey@356 mAd137_1 mAd137_2 d1 e2 basic__key adr=137
Xkey@357 mAd136_1 mAd136_2 d3 e2 basic__key adr=136
Xkey@358 mAd130_1 mAd130_2 a3 e4 basic__key adr=130
Xkey@359 mAd247_1 mAd247_2 a5 e4 basic__key adr=247
Xkey@360 mAd241_1 mAd241_2 d5 e6 basic__key adr=241
Xkey@361 mAd240_1 mAd240_2 d7 e6 basic__key adr=240
Xkey@362 mAd351_1 mAd351_2 a7 Z5 basic__key adr=351
Xkey@363 mAd340_1 mAd340_2 K13 Z5 basic__key adr=340
Xkey@364 mAd320_1 mAd320_2 K13 Z6 basic__key adr=320
Xkey@365 mAd337_1 mAd337_2 e7 f6 basic__key adr=337
Xkey@366 mAd220_1 mAd220_2 d7 f6 basic__key adr=220
Xkey@367 mAd221_1 mAd221_2 d5 f6 basic__key adr=221
Xkey@368 mAd222_1 mAd222_2 e5 f6 basic__key adr=222
Xkey@369 mAd155_1 mAd155_2 e3 f2 basic__key adr=155
Xkey@370 mAd156_1 mAd156_2 d3 f2 basic__key adr=156
Xkey@371 mAd157_1 mAd157_2 d1 f2 basic__key adr=157
Xkey@372 mAd040_1 mAd040_2 e1 f2 basic__key adr=40
Xkey@373 mAd440_1 mAd440_2 e1 g2 basic__key adr=440
Xkey@374 mAd557_1 mAd557_2 d1 g2 basic__key adr=557
Xkey@375 mAd556_1 mAd556_2 d3 g2 basic__key adr=556
Xkey@376 mAd555_1 mAd555_2 e3 g2 basic__key adr=555
Xkey@377 mAd622_1 mAd622_2 e5 g6 basic__key adr=622
Xkey@378 mAd621_1 mAd621_2 d5 g6 basic__key adr=621
Xkey@379 mAd620_1 mAd620_2 d7 g6 basic__key adr=620
Xkey@380 mAd737_1 mAd737_2 e7 g6 basic__key adr=737
Xkey@381 mAd720_1 mAd720_2 K13 Z7 basic__key adr=720
Xkey@382 mAd426_1 mAd426_2 g1 X8 basic__key adr=426
Xkey@383 mAd537_1 mAd537_2 d1 h2 basic__key adr=537
Xkey@384 mAd536_1 mAd536_2 d3 h2 basic__key adr=536
Xkey@385 mAd530_1 mAd530_2 g3 h4 basic__key adr=530
Xkey@386 mAd647_1 mAd647_2 g5 h4 basic__key adr=647
Xkey@387 mAd641_1 mAd641_2 d5 h6 basic__key adr=641
Xkey@388 mAd640_1 mAd640_2 d7 h6 basic__key adr=640
Xkey@389 mAd751_1 mAd751_2 g7 Z8 basic__key adr=751
Xkey@390 mAd740_1 mAd740_2 K13 Z8 basic__key adr=740
Xkey@391 mAd406_1 mAd406_2 g1 X9 basic__key adr=406
Xkey@392 mAd405_1 mAd405_2 h1 X9 basic__key adr=405
Xkey@393 mAd531_1 mAd531_2 h3 i4 basic__key adr=531
Xkey@394 mAd508_1 mAd508_2 g3 i4 basic__key adr=508
Xkey@395 mAd667_1 mAd667_2 g5 i4 basic__key adr=667
Xkey@396 mAd646_1 mAd646_2 h5 i4 basic__key adr=646
Xkey@397 mAd772_1 mAd772_2 h7 Z9 basic__key adr=772
Xkey@398 mAd771_1 mAd771_2 g7 Z9 basic__key adr=771
Xkey@399 mAd760_1 mAd760_2 K13 Z9 basic__key adr=760
Xkey@400 mAd416_1 mAd416_2 g1 X10 basic__key adr=416
Xkey@401 mAd415_1 mAd415_2 h1 X10 basic__key adr=415
Xkey@402 mAd541_1 mAd541_2 h3 j2 basic__key adr=541
Xkey@403 mAd520_1 mAd520_2 g3 j2 basic__key adr=520
Xkey@404 mAd657_1 mAd657_2 g5 j2 basic__key adr=657
Xkey@405 mAd636_1 mAd636_2 h5 j2 basic__key adr=636
Xkey@406 mAd762_1 mAd762_2 h7 Z10 basic__key adr=762
Xkey@407 mAd761_1 mAd761_2 g7 Z10 basic__key adr=761
Xkey@408 mAd750_1 mAd750_2 K13 Z10 basic__key adr=750
Xkey@409 mAd730_1 mAd730_2 K13 Z11 basic__key adr=730
Xkey@410 mAd741_1 mAd741_2 g7 Z11 basic__key adr=741
Xkey@411 mAd630_1 mAd630_2 K10 k3 basic__key adr=630
Xkey@412 mAd631_1 mAd631_2 K9 k3 basic__key adr=631
Xkey@413 mAd637_1 mAd637_2 g5 k2 basic__key adr=637
Xkey@414 mAd540_1 mAd540_2 g3 k2 basic__key adr=540
Xkey@415 mAd546_1 mAd546_2 K4 k1 basic__key adr=546
Xkey@416 mAd547_1 mAd547_2 K3 k1 basic__key adr=547
Xkey@417 mAd436_1 mAd436_2 g1 X11 basic__key adr=436
Xkey@418 mAd450_1 mAd450_2 K2 l1 basic__key adr=450
Xkey@419 mAd567_1 mAd567_2 K3 l1 basic__key adr=567
Xkey@420 mAd566_1 mAd566_2 K4 l1 basic__key adr=566
Xkey@421 mAd565_1 mAd565_2 K5 l1 basic__key adr=565
Xkey@422 mAd612_1 mAd612_2 K8 l3 basic__key adr=612
Xkey@423 mAd611_1 mAd611_2 K9 l3 basic__key adr=611
Xkey@424 mAd610_1 mAd610_2 K10 l3 basic__key adr=610
Xkey@425 mAd727_1 mAd727_2 K11 l3 basic__key adr=727
Xkey@426 mAd710_1 mAd710_2 K13 Z12 basic__key adr=710
Xkey@427 mAd700_1 mAd700_2 K13 X13 basic__key adr=700
Xkey@428 mAd711_1 mAd711_2 K12 X13 basic__key adr=711
Xkey@429 mAd717_1 mAd717_2 K11 X13 basic__key adr=717
Xkey@430 mAd600_1 mAd600_2 K10 X13 basic__key adr=600
Xkey@431 mAd601_1 mAd601_2 K9 X13 basic__key adr=601
Xkey@432 mAd602_1 mAd602_2 K8 X13 basic__key adr=602
Xkey@433 mAd607_1 mAd607_2 K7 X13 basic__key adr=607
Xkey@434 mAd570_1 mAd570_2 K6 X13 basic__key adr=570
Xkey@435 mAd575_1 mAd575_2 K5 X13 basic__key adr=575
Xkey@436 mAd576_1 mAd576_2 K4 X13 basic__key adr=576
Xkey@437 mAd577_1 mAd577_2 K3 X13 basic__key adr=577
Xkey@438 mAd460_1 mAd460_2 K2 X13 basic__key adr=460
Xkey@439 mAd466_1 mAd466_2 K1 X13 basic__key adr=466
.ENDS _5400TP094__CB

.global gnd

*** TOP LEVEL CELL: 5400TP094NEW{sch}
.options filetype=ascii
.tran 0.1u 4u
.include "C:/IvanovFolder/PADIC/Spice64/models/soimod018.tec"
.global VDDA! VSSA!
.options method=gear reltol=0.01 itl4=500 altinit=10 RSHUNT=1.41G cshunt=1e-15 abstol=5u chgtol=2p vntol=5u trtol=7
XCB@0 CB@0_K0 CB@0_K1 CB@0_K10 CB@0_K11 CB@0_K12 CB@0_K13 CB@0_K2 CB@0_K3 CB@0_K4 CB@0_K5 CB@0_K6 CB@0_K7 CB@0_K8 CB@0_K9 CB@0_mAd000_1 CB@0_mAd000_2 CB@0_mAd001_1 CB@0_mAd001_2 CB@0_mAd002_1 CB@0_mAd002_2 CB@0_mAd003_1 CB@0_mAd003_2 CB@0_mAd004_1 CB@0_mAd004_2 CB@0_mAd005_1 CB@0_mAd005_2 CB@0_mAd006_1 CB@0_mAd006_2 CB@0_mAd007_1 CB@0_mAd007_2 CB@0_mAd010_1 CB@0_mAd010_2 CB@0_mAd011_1 CB@0_mAd011_2 CB@0_mAd012_1 CB@0_mAd012_2 CB@0_mAd013_1 CB@0_mAd013_2 CB@0_mAd014_1 CB@0_mAd014_2 CB@0_mAd015_1 
+CB@0_mAd015_2 CB@0_mAd016_1 CB@0_mAd016_2 CB@0_mAd017_1 CB@0_mAd017_2 CB@0_mAd020_1 CB@0_mAd020_2 CB@0_mAd021_1 CB@0_mAd021_2 CB@0_mAd022_1 CB@0_mAd022_2 CB@0_mAd023_1 CB@0_mAd023_2 CB@0_mAd024_1 CB@0_mAd024_2 CB@0_mAd025_1 CB@0_mAd025_2 CB@0_mAd026_1 CB@0_mAd026_2 CB@0_mAd027_1 CB@0_mAd027_2 CB@0_mAd030_1 CB@0_mAd030_2 CB@0_mAd031_1 CB@0_mAd031_2 CB@0_mAd032_1 CB@0_mAd032_2 CB@0_mAd033_1 CB@0_mAd033_2 CB@0_mAd034_1 CB@0_mAd034_2 CB@0_mAd035_1 CB@0_mAd035_2 CB@0_mAd036_1 CB@0_mAd036_2 CB@0_mAd037_1 
+CB@0_mAd037_2 CB@0_mAd040_1 CB@0_mAd040_2 CB@0_mAd041_1 CB@0_mAd041_2 CB@0_mAd042_1 CB@0_mAd042_2 CB@0_mAd043_1 CB@0_mAd043_2 CB@0_mAd044_1 CB@0_mAd044_2 CB@0_mAd045_1 CB@0_mAd045_2 CB@0_mAd046_1 CB@0_mAd046_2 CB@0_mAd047_1 CB@0_mAd047_2 CB@0_mAd050_1 CB@0_mAd050_2 CB@0_mAd051_1 CB@0_mAd051_2 CB@0_mAd052_1 CB@0_mAd052_2 CB@0_mAd053_1 CB@0_mAd053_2 CB@0_mAd054_1 CB@0_mAd054_2 net@1451 net@1451 CB@0_mAd056_1 CB@0_mAd056_2 CB@0_mAd057_1 CB@0_mAd057_2 CB@0_mAd060_1 CB@0_mAd060_2 CB@0_mAd066_1 CB@0_mAd066_2 
+CB@0_mAd067_1 CB@0_mAd067_2 net@1452 net@1452 CB@0_mAd101_1 CB@0_mAd101_2 CB@0_mAd102_1 CB@0_mAd102_2 CB@0_mAd110_1 CB@0_mAd110_2 CB@0_mAd111_1 CB@0_mAd111_2 CB@0_mAd112_1 CB@0_mAd112_2 CB@0_mAd113_1 CB@0_mAd113_2 CB@0_mAd114_1 CB@0_mAd114_2 CB@0_mAd115_1 CB@0_mAd115_2 CB@0_mAd116_1 CB@0_mAd116_2 CB@0_mAd117_1 CB@0_mAd117_2 CB@0_mAd120_1 CB@0_mAd120_2 CB@0_mAd121_1 CB@0_mAd121_2 CB@0_mAd122_1 CB@0_mAd122_2 CB@0_mAd123_1 CB@0_mAd123_2 CB@0_mAd124_1 CB@0_mAd124_2 CB@0_mAd125_1 CB@0_mAd125_2 CB@0_mAd126_1 
+CB@0_mAd126_2 CB@0_mAd127_1 CB@0_mAd127_2 CB@0_mAd130_1 CB@0_mAd130_2 CB@0_mAd131_1 CB@0_mAd131_2 CB@0_mAd132_1 CB@0_mAd132_2 CB@0_mAd133_1 CB@0_mAd133_2 CB@0_mAd134_1 CB@0_mAd134_2 CB@0_mAd135_1 CB@0_mAd135_2 CB@0_mAd136_1 CB@0_mAd136_2 CB@0_mAd137_1 CB@0_mAd137_2 CB@0_mAd140_1 CB@0_mAd140_2 CB@0_mAd141_1 CB@0_mAd141_2 CB@0_mAd142_1 CB@0_mAd142_2 CB@0_mAd143_1 CB@0_mAd143_2 CB@0_mAd144_1 CB@0_mAd144_2 CB@0_mAd145_1 CB@0_mAd145_2 CB@0_mAd146_1 CB@0_mAd146_2 CB@0_mAd147_1 CB@0_mAd147_2 CB@0_mAd150_1 
+CB@0_mAd150_2 CB@0_mAd151_1 CB@0_mAd151_2 CB@0_mAd152_1 CB@0_mAd152_2 CB@0_mAd153_1 CB@0_mAd153_2 CB@0_mAd154_1 CB@0_mAd154_2 CB@0_mAd155_1 CB@0_mAd155_2 CB@0_mAd156_1 CB@0_mAd156_2 CB@0_mAd157_1 CB@0_mAd157_2 CB@0_mAd160_1 CB@0_mAd160_2 CB@0_mAd161_1 CB@0_mAd161_2 CB@0_mAd162_1 CB@0_mAd162_2 CB@0_mAd163_1 CB@0_mAd163_2 CB@0_mAd164_1 CB@0_mAd164_2 CB@0_mAd165_1 CB@0_mAd165_2 CB@0_mAd166_1 CB@0_mAd166_2 CB@0_mAd167_1 CB@0_mAd167_2 CB@0_mAd170_1 CB@0_mAd170_2 CB@0_mAd171_1 CB@0_mAd171_2 CB@0_mAd172_1 
+CB@0_mAd172_2 CB@0_mAd173_1 CB@0_mAd173_2 CB@0_mAd175_1 CB@0_mAd175_2 CB@0_mAd176_1 CB@0_mAd176_2 CB@0_mAd177_1 CB@0_mAd177_2 CB@0_mAd200_1 CB@0_mAd200_2 CB@0_mAd201_1 CB@0_mAd201_2 CB@0_mAd202_1 CB@0_mAd202_2 CB@0_mAd204_1 CB@0_mAd204_2 CB@0_mAd205_1 CB@0_mAd205_2 CB@0_mAd206_1 CB@0_mAd206_2 CB@0_mAd207_1 CB@0_mAd207_2 CB@0_mAd210_1 CB@0_mAd210_2 CB@0_mAd211_1 CB@0_mAd211_2 CB@0_mAd212_1 CB@0_mAd212_2 CB@0_mAd213_1 CB@0_mAd213_2 CB@0_mAd214_1 CB@0_mAd214_2 CB@0_mAd215_1 CB@0_mAd215_2 CB@0_mAd216_1 
+CB@0_mAd216_2 CB@0_mAd217_1 CB@0_mAd217_2 CB@0_mAd220_1 CB@0_mAd220_2 CB@0_mAd221_1 CB@0_mAd221_2 CB@0_mAd222_1 CB@0_mAd222_2 CB@0_mAd223_1 CB@0_mAd223_2 CB@0_mAd224_1 CB@0_mAd224_2 CB@0_mAd225_1 CB@0_mAd225_2 CB@0_mAd226_1 CB@0_mAd226_2 CB@0_mAd227_1 CB@0_mAd227_2 CB@0_mAd230_1 CB@0_mAd230_2 CB@0_mAd231_1 CB@0_mAd231_2 CB@0_mAd232_1 CB@0_mAd232_2 CB@0_mAd233_1 CB@0_mAd233_2 CB@0_mAd234_1 CB@0_mAd234_2 CB@0_mAd235_1 CB@0_mAd235_2 CB@0_mAd236_1 CB@0_mAd236_2 CB@0_mAd237_1 CB@0_mAd237_2 CB@0_mAd240_1 
+CB@0_mAd240_2 CB@0_mAd241_1 CB@0_mAd241_2 CB@0_mAd242_1 CB@0_mAd242_2 CB@0_mAd243_1 CB@0_mAd243_2 CB@0_mAd244_1 CB@0_mAd244_2 CB@0_mAd245_1 CB@0_mAd245_2 CB@0_mAd246_1 CB@0_mAd246_2 CB@0_mAd247_1 CB@0_mAd247_2 CB@0_mAd250_1 CB@0_mAd250_2 CB@0_mAd251_1 CB@0_mAd251_2 CB@0_mAd252_1 CB@0_mAd252_2 CB@0_mAd253_1 CB@0_mAd253_2 CB@0_mAd254_1 CB@0_mAd254_2 CB@0_mAd255_1 CB@0_mAd255_2 CB@0_mAd256_1 CB@0_mAd256_2 CB@0_mAd257_1 CB@0_mAd257_2 CB@0_mAd260_1 CB@0_mAd260_2 CB@0_mAd261_1 CB@0_mAd261_2 CB@0_mAd262_1 
+CB@0_mAd262_2 CB@0_mAd263_1 CB@0_mAd263_2 CB@0_mAd264_1 CB@0_mAd264_2 CB@0_mAd265_1 CB@0_mAd265_2 CB@0_mAd266_1 CB@0_mAd266_2 CB@0_mAd267_1 CB@0_mAd267_2 CB@0_mAd275_1 CB@0_mAd275_2 CB@0_mAd276_1 CB@0_mAd276_2 net@1453 net@1453 net@1456 net@1456 net@1455 net@1455 CB@0_mAd311_1 CB@0_mAd311_2 CB@0_mAd317_1 CB@0_mAd317_2 CB@0_mAd320_1 CB@0_mAd320_2 CB@0_mAd321_1 CB@0_mAd321_2 net@1454 net@1454 CB@0_mAd323_1 CB@0_mAd323_2 CB@0_mAd324_1 CB@0_mAd324_2 CB@0_mAd325_1 CB@0_mAd325_2 CB@0_mAd326_1 CB@0_mAd326_2 
+CB@0_mAd327_1 CB@0_mAd327_2 CB@0_mAd330_1 CB@0_mAd330_2 CB@0_mAd331_1 CB@0_mAd331_2 CB@0_mAd332_1 CB@0_mAd332_2 CB@0_mAd333_1 CB@0_mAd333_2 CB@0_mAd334_1 CB@0_mAd334_2 CB@0_mAd335_1 CB@0_mAd335_2 CB@0_mAd336_1 CB@0_mAd336_2 CB@0_mAd337_1 CB@0_mAd337_2 CB@0_mAd340_1 CB@0_mAd340_2 CB@0_mAd341_1 CB@0_mAd341_2 CB@0_mAd342_1 CB@0_mAd342_2 CB@0_mAd343_1 CB@0_mAd343_2 CB@0_mAd344_1 CB@0_mAd344_2 CB@0_mAd345_1 CB@0_mAd345_2 CB@0_mAd346_1 CB@0_mAd346_2 CB@0_mAd347_1 CB@0_mAd347_2 CB@0_mAd350_1 CB@0_mAd350_2 
+CB@0_mAd351_1 CB@0_mAd351_2 CB@0_mAd352_1 CB@0_mAd352_2 CB@0_mAd353_1 CB@0_mAd353_2 CB@0_mAd354_1 CB@0_mAd354_2 CB@0_mAd355_1 CB@0_mAd355_2 CB@0_mAd356_1 CB@0_mAd356_2 CB@0_mAd357_1 CB@0_mAd357_2 CB@0_mAd360_1 CB@0_mAd360_2 CB@0_mAd361_1 CB@0_mAd361_2 CB@0_mAd362_1 CB@0_mAd362_2 CB@0_mAd363_1 CB@0_mAd363_2 CB@0_mAd364_1 CB@0_mAd364_2 CB@0_mAd365_1 CB@0_mAd365_2 CB@0_mAd366_1 CB@0_mAd366_2 CB@0_mAd367_1 CB@0_mAd367_2 CB@0_mAd371_1 CB@0_mAd371_2 CB@0_mAd372_1 CB@0_mAd372_2 CB@0_mAd373_1 CB@0_mAd373_2 
+CB@0_mAd374_1 CB@0_mAd374_2 CB@0_mAd375_1 CB@0_mAd375_2 CB@0_mAd376_1 CB@0_mAd376_2 CB@0_mAd377_1 CB@0_mAd377_2 CB@0_mAd400_1 CB@0_mAd400_2 CB@0_mAd401_1 CB@0_mAd401_2 CB@0_mAd402_1 CB@0_mAd402_2 CB@0_mAd403_1 CB@0_mAd403_2 CB@0_mAd404_1 CB@0_mAd404_2 CB@0_mAd405_1 CB@0_mAd405_2 CB@0_mAd406_1 CB@0_mAd406_2 CB@0_mAd407_1 CB@0_mAd407_2 CB@0_mAd410_1 CB@0_mAd410_2 CB@0_mAd411_1 CB@0_mAd411_2 CB@0_mAd412_1 CB@0_mAd412_2 CB@0_mAd413_1 CB@0_mAd413_2 CB@0_mAd414_1 CB@0_mAd414_2 CB@0_mAd415_1 CB@0_mAd415_2 
+CB@0_mAd416_1 CB@0_mAd416_2 CB@0_mAd417_1 CB@0_mAd417_2 CB@0_mAd420_1 CB@0_mAd420_2 CB@0_mAd421_1 CB@0_mAd421_2 CB@0_mAd422_1 CB@0_mAd422_2 CB@0_mAd423_1 CB@0_mAd423_2 CB@0_mAd424_1 CB@0_mAd424_2 CB@0_mAd425_1 CB@0_mAd425_2 CB@0_mAd426_1 CB@0_mAd426_2 CB@0_mAd427_1 CB@0_mAd427_2 CB@0_mAd430_1 CB@0_mAd430_2 CB@0_mAd431_1 CB@0_mAd431_2 CB@0_mAd432_1 CB@0_mAd432_2 CB@0_mAd433_1 CB@0_mAd433_2 CB@0_mAd434_1 CB@0_mAd434_2 CB@0_mAd435_1 CB@0_mAd435_2 CB@0_mAd436_1 CB@0_mAd436_2 CB@0_mAd437_1 CB@0_mAd437_2 
+CB@0_mAd440_1 CB@0_mAd440_2 CB@0_mAd441_1 CB@0_mAd441_2 CB@0_mAd442_1 CB@0_mAd442_2 CB@0_mAd443_1 CB@0_mAd443_2 CB@0_mAd444_1 CB@0_mAd444_2 CB@0_mAd445_1 CB@0_mAd445_2 CB@0_mAd446_1 CB@0_mAd446_2 CB@0_mAd447_1 CB@0_mAd447_2 CB@0_mAd450_1 CB@0_mAd450_2 CB@0_mAd451_1 CB@0_mAd451_2 CB@0_mAd452_1 CB@0_mAd452_2 CB@0_mAd453_1 CB@0_mAd453_2 CB@0_mAd454_1 CB@0_mAd454_2 CB@0_mAd455_1 CB@0_mAd455_2 CB@0_mAd456_1 CB@0_mAd456_2 CB@0_mAd457_1 CB@0_mAd457_2 CB@0_mAd460_1 CB@0_mAd460_2 CB@0_mAd466_1 CB@0_mAd466_2 
+CB@0_mAd467_1 CB@0_mAd467_2 CB@0_mAd500_1 CB@0_mAd500_2 CB@0_mAd501_1 CB@0_mAd501_2 CB@0_mAd502_1 CB@0_mAd502_2 CB@0_mAd508_1 CB@0_mAd508_2 CB@0_mAd509_1 CB@0_mAd509_2 CB@0_mAd512_1 CB@0_mAd512_2 CB@0_mAd513_1 CB@0_mAd513_2 CB@0_mAd514_1 CB@0_mAd514_2 CB@0_mAd515_1 CB@0_mAd515_2 CB@0_mAd516_1 CB@0_mAd516_2 CB@0_mAd517_1 CB@0_mAd517_2 CB@0_mAd520_1 CB@0_mAd520_2 CB@0_mAd521_1 CB@0_mAd521_2 CB@0_mAd522_1 CB@0_mAd522_2 CB@0_mAd523_1 CB@0_mAd523_2 CB@0_mAd524_1 CB@0_mAd524_2 CB@0_mAd525_1 CB@0_mAd525_2 
+CB@0_mAd526_1 CB@0_mAd526_2 CB@0_mAd527_1 CB@0_mAd527_2 CB@0_mAd530_1 CB@0_mAd530_2 CB@0_mAd531_1 CB@0_mAd531_2 CB@0_mAd532_1 CB@0_mAd532_2 CB@0_mAd533_1 CB@0_mAd533_2 CB@0_mAd534_1 CB@0_mAd534_2 CB@0_mAd535_1 CB@0_mAd535_2 CB@0_mAd536_1 CB@0_mAd536_2 CB@0_mAd537_1 CB@0_mAd537_2 CB@0_mAd540_1 CB@0_mAd540_2 CB@0_mAd541_1 CB@0_mAd541_2 CB@0_mAd542_1 CB@0_mAd542_2 CB@0_mAd543_1 CB@0_mAd543_2 CB@0_mAd544_1 CB@0_mAd544_2 CB@0_mAd545_1 CB@0_mAd545_2 CB@0_mAd546_1 CB@0_mAd546_2 CB@0_mAd547_1 CB@0_mAd547_2 
+CB@0_mAd550_1 CB@0_mAd550_2 CB@0_mAd551_1 CB@0_mAd551_2 CB@0_mAd552_1 CB@0_mAd552_2 CB@0_mAd553_1 CB@0_mAd553_2 CB@0_mAd554_1 CB@0_mAd554_2 CB@0_mAd555_1 CB@0_mAd555_2 CB@0_mAd556_1 CB@0_mAd556_2 CB@0_mAd557_1 CB@0_mAd557_2 CB@0_mAd560_1 CB@0_mAd560_2 CB@0_mAd561_1 CB@0_mAd561_2 CB@0_mAd562_1 CB@0_mAd562_2 CB@0_mAd563_1 CB@0_mAd563_2 CB@0_mAd564_1 CB@0_mAd564_2 CB@0_mAd565_1 CB@0_mAd565_2 CB@0_mAd566_1 CB@0_mAd566_2 CB@0_mAd567_1 CB@0_mAd567_2 CB@0_mAd570_1 CB@0_mAd570_2 CB@0_mAd571_1 CB@0_mAd571_2 
+CB@0_mAd572_1 CB@0_mAd572_2 CB@0_mAd573_1 CB@0_mAd573_2 CB@0_mAd575_1 CB@0_mAd575_2 CB@0_mAd576_1 CB@0_mAd576_2 CB@0_mAd577_1 CB@0_mAd577_2 CB@0_mAd600_1 CB@0_mAd600_2 CB@0_mAd601_1 CB@0_mAd601_2 CB@0_mAd602_1 CB@0_mAd602_2 CB@0_mAd604_1 CB@0_mAd604_2 CB@0_mAd605_1 CB@0_mAd605_2 CB@0_mAd606_1 CB@0_mAd606_2 CB@0_mAd607_1 CB@0_mAd607_2 CB@0_mAd610_1 CB@0_mAd610_2 CB@0_mAd611_1 CB@0_mAd611_2 CB@0_mAd612_1 CB@0_mAd612_2 CB@0_mAd613_1 CB@0_mAd613_2 CB@0_mAd614_1 CB@0_mAd614_2 CB@0_mAd615_1 CB@0_mAd615_2 
+CB@0_mAd616_1 CB@0_mAd616_2 CB@0_mAd617_1 CB@0_mAd617_2 CB@0_mAd620_1 CB@0_mAd620_2 CB@0_mAd621_1 CB@0_mAd621_2 CB@0_mAd622_1 CB@0_mAd622_2 CB@0_mAd623_1 CB@0_mAd623_2 CB@0_mAd624_1 CB@0_mAd624_2 CB@0_mAd625_1 CB@0_mAd625_2 CB@0_mAd626_1 CB@0_mAd626_2 CB@0_mAd627_1 CB@0_mAd627_2 CB@0_mAd630_1 CB@0_mAd630_2 CB@0_mAd631_1 CB@0_mAd631_2 CB@0_mAd632_1 CB@0_mAd632_2 CB@0_mAd633_1 CB@0_mAd633_2 CB@0_mAd634_1 CB@0_mAd634_2 CB@0_mAd635_1 CB@0_mAd635_2 CB@0_mAd636_1 CB@0_mAd636_2 CB@0_mAd637_1 CB@0_mAd637_2 
+CB@0_mAd640_1 CB@0_mAd640_2 CB@0_mAd641_1 CB@0_mAd641_2 CB@0_mAd642_1 CB@0_mAd642_2 CB@0_mAd643_1 CB@0_mAd643_2 CB@0_mAd644_1 CB@0_mAd644_2 CB@0_mAd645_1 CB@0_mAd645_2 CB@0_mAd646_1 CB@0_mAd646_2 CB@0_mAd647_1 CB@0_mAd647_2 CB@0_mAd650_1 CB@0_mAd650_2 CB@0_mAd651_1 CB@0_mAd651_2 CB@0_mAd652_1 CB@0_mAd652_2 CB@0_mAd653_1 CB@0_mAd653_2 CB@0_mAd654_1 CB@0_mAd654_2 CB@0_mAd655_1 CB@0_mAd655_2 CB@0_mAd656_1 CB@0_mAd656_2 CB@0_mAd657_1 CB@0_mAd657_2 CB@0_mAd660_1 CB@0_mAd660_2 CB@0_mAd661_1 CB@0_mAd661_2 
+CB@0_mAd662_1 CB@0_mAd662_2 CB@0_mAd663_1 CB@0_mAd663_2 CB@0_mAd664_1 CB@0_mAd664_2 CB@0_mAd665_1 CB@0_mAd665_2 CB@0_mAd666_1 CB@0_mAd666_2 CB@0_mAd667_1 CB@0_mAd667_2 CB@0_mAd675_1 CB@0_mAd675_2 CB@0_mAd676_1 CB@0_mAd676_2 CB@0_mAd677_1 CB@0_mAd677_2 CB@0_mAd700_1 CB@0_mAd700_2 CB@0_mAd710_1 CB@0_mAd710_2 CB@0_mAd711_1 CB@0_mAd711_2 CB@0_mAd717_1 CB@0_mAd717_2 CB@0_mAd720_1 CB@0_mAd720_2 CB@0_mAd721_1 CB@0_mAd721_2 CB@0_mAd722_1 CB@0_mAd722_2 CB@0_mAd723_1 CB@0_mAd723_2 CB@0_mAd724_1 CB@0_mAd724_2 
+CB@0_mAd725_1 CB@0_mAd725_2 CB@0_mAd726_1 CB@0_mAd726_2 CB@0_mAd727_1 CB@0_mAd727_2 CB@0_mAd730_1 CB@0_mAd730_2 CB@0_mAd731_1 CB@0_mAd731_2 CB@0_mAd732_1 CB@0_mAd732_2 CB@0_mAd733_1 CB@0_mAd733_2 CB@0_mAd734_1 CB@0_mAd734_2 CB@0_mAd735_1 CB@0_mAd735_2 CB@0_mAd736_1 CB@0_mAd736_2 CB@0_mAd737_1 CB@0_mAd737_2 CB@0_mAd740_1 CB@0_mAd740_2 CB@0_mAd741_1 CB@0_mAd741_2 CB@0_mAd742_1 CB@0_mAd742_2 CB@0_mAd743_1 CB@0_mAd743_2 CB@0_mAd744_1 CB@0_mAd744_2 CB@0_mAd745_1 CB@0_mAd745_2 CB@0_mAd746_1 CB@0_mAd746_2 
+CB@0_mAd747_1 CB@0_mAd747_2 CB@0_mAd750_1 CB@0_mAd750_2 CB@0_mAd751_1 CB@0_mAd751_2 CB@0_mAd752_1 CB@0_mAd752_2 CB@0_mAd753_1 CB@0_mAd753_2 CB@0_mAd754_1 CB@0_mAd754_2 CB@0_mAd755_1 CB@0_mAd755_2 CB@0_mAd756_1 CB@0_mAd756_2 CB@0_mAd757_1 CB@0_mAd757_2 CB@0_mAd760_1 CB@0_mAd760_2 CB@0_mAd761_1 CB@0_mAd761_2 CB@0_mAd762_1 CB@0_mAd762_2 CB@0_mAd763_1 CB@0_mAd763_2 CB@0_mAd764_1 CB@0_mAd764_2 CB@0_mAd765_1 CB@0_mAd765_2 CB@0_mAd766_1 CB@0_mAd766_2 CB@0_mAd767_1 CB@0_mAd767_2 CB@0_mAd771_1 CB@0_mAd771_2 
+CB@0_mAd772_1 CB@0_mAd772_2 CB@0_mAd773_1 CB@0_mAd773_2 CB@0_mAd774_1 CB@0_mAd774_2 CB@0_mAd775_1 CB@0_mAd775_2 CB@0_mAd776_1 CB@0_mAd776_2 CB@0_mAd777_1 CB@0_mAd777_2 net@1447 in1 CB@0_X10 CB@0_X11 CB@0_X12 CB@0_X13 CB@0_X2 CB@0_X3 CB@0_X4 CB@0_X5 CB@0_X6 CB@0_X7 CB@0_X8 CB@0_X9 CB@0_Y1 CB@0_Y10 CB@0_Y11 CB@0_Y12 CB@0_Y2 CB@0_Y3 CB@0_Y4 CB@0_Y5 CB@0_Y6 CB@0_Y7 CB@0_Y8 CB@0_Y9 CB@0_Z1 CB@0_Z10 CB@0_Z11 CB@0_Z12 CB@0_Z2 CB@0_Z3 CB@0_Z4 CB@0_Z5 CB@0_Z6 CB@0_Z7 CB@0_Z8 CB@0_Z9 _5400TP094__CB
XCB@1 CB@1_K0 CB@1_K1 CB@1_K10 CB@1_K11 CB@1_K12 CB@1_K13 CB@1_K2 CB@1_K3 CB@1_K4 CB@1_K5 CB@1_K6 CB@1_K7 CB@1_K8 CB@1_K9 CB@1_mAd000_1 CB@1_mAd000_2 CB@1_mAd001_1 CB@1_mAd001_2 CB@1_mAd002_1 CB@1_mAd002_2 CB@1_mAd003_1 CB@1_mAd003_2 CB@1_mAd004_1 CB@1_mAd004_2 CB@1_mAd005_1 CB@1_mAd005_2 CB@1_mAd006_1 CB@1_mAd006_2 CB@1_mAd007_1 CB@1_mAd007_2 CB@1_mAd010_1 CB@1_mAd010_2 CB@1_mAd011_1 CB@1_mAd011_2 CB@1_mAd012_1 CB@1_mAd012_2 net@1457 net@1457 CB@1_mAd014_1 CB@1_mAd014_2 CB@1_mAd015_1 CB@1_mAd015_2 
+CB@1_mAd016_1 CB@1_mAd016_2 CB@1_mAd017_1 CB@1_mAd017_2 CB@1_mAd020_1 CB@1_mAd020_2 CB@1_mAd021_1 CB@1_mAd021_2 CB@1_mAd022_1 CB@1_mAd022_2 CB@1_mAd023_1 CB@1_mAd023_2 CB@1_mAd024_1 CB@1_mAd024_2 CB@1_mAd025_1 CB@1_mAd025_2 CB@1_mAd026_1 CB@1_mAd026_2 CB@1_mAd027_1 CB@1_mAd027_2 CB@1_mAd030_1 CB@1_mAd030_2 CB@1_mAd031_1 CB@1_mAd031_2 CB@1_mAd032_1 CB@1_mAd032_2 CB@1_mAd033_1 CB@1_mAd033_2 CB@1_mAd034_1 CB@1_mAd034_2 CB@1_mAd035_1 CB@1_mAd035_2 CB@1_mAd036_1 CB@1_mAd036_2 CB@1_mAd037_1 CB@1_mAd037_2 
+CB@1_mAd040_1 CB@1_mAd040_2 CB@1_mAd041_1 CB@1_mAd041_2 CB@1_mAd042_1 CB@1_mAd042_2 CB@1_mAd043_1 CB@1_mAd043_2 CB@1_mAd044_1 CB@1_mAd044_2 CB@1_mAd045_1 CB@1_mAd045_2 CB@1_mAd046_1 CB@1_mAd046_2 CB@1_mAd047_1 CB@1_mAd047_2 CB@1_mAd050_1 CB@1_mAd050_2 CB@1_mAd051_1 CB@1_mAd051_2 CB@1_mAd052_1 CB@1_mAd052_2 CB@1_mAd053_1 CB@1_mAd053_2 CB@1_mAd054_1 CB@1_mAd054_2 CB@1_mAd055_1 CB@1_mAd055_2 CB@1_mAd056_1 CB@1_mAd056_2 CB@1_mAd057_1 CB@1_mAd057_2 CB@1_mAd060_1 CB@1_mAd060_2 CB@1_mAd066_1 CB@1_mAd066_2 
+CB@1_mAd067_1 CB@1_mAd067_2 CB@1_mAd100_1 CB@1_mAd100_2 CB@1_mAd101_1 CB@1_mAd101_2 net@1458 net@1458 CB@1_mAd110_1 CB@1_mAd110_2 CB@1_mAd111_1 CB@1_mAd111_2 CB@1_mAd112_1 CB@1_mAd112_2 CB@1_mAd113_1 CB@1_mAd113_2 CB@1_mAd114_1 CB@1_mAd114_2 CB@1_mAd115_1 CB@1_mAd115_2 CB@1_mAd116_1 CB@1_mAd116_2 CB@1_mAd117_1 CB@1_mAd117_2 CB@1_mAd120_1 CB@1_mAd120_2 CB@1_mAd121_1 CB@1_mAd121_2 CB@1_mAd122_1 CB@1_mAd122_2 CB@1_mAd123_1 CB@1_mAd123_2 CB@1_mAd124_1 CB@1_mAd124_2 CB@1_mAd125_1 CB@1_mAd125_2 CB@1_mAd126_1 
+CB@1_mAd126_2 CB@1_mAd127_1 CB@1_mAd127_2 CB@1_mAd130_1 CB@1_mAd130_2 CB@1_mAd131_1 CB@1_mAd131_2 CB@1_mAd132_1 CB@1_mAd132_2 CB@1_mAd133_1 CB@1_mAd133_2 CB@1_mAd134_1 CB@1_mAd134_2 CB@1_mAd135_1 CB@1_mAd135_2 CB@1_mAd136_1 CB@1_mAd136_2 CB@1_mAd137_1 CB@1_mAd137_2 CB@1_mAd140_1 CB@1_mAd140_2 CB@1_mAd141_1 CB@1_mAd141_2 CB@1_mAd142_1 CB@1_mAd142_2 CB@1_mAd143_1 CB@1_mAd143_2 CB@1_mAd144_1 CB@1_mAd144_2 CB@1_mAd145_1 CB@1_mAd145_2 CB@1_mAd146_1 CB@1_mAd146_2 CB@1_mAd147_1 CB@1_mAd147_2 CB@1_mAd150_1 
+CB@1_mAd150_2 CB@1_mAd151_1 CB@1_mAd151_2 CB@1_mAd152_1 CB@1_mAd152_2 CB@1_mAd153_1 CB@1_mAd153_2 CB@1_mAd154_1 CB@1_mAd154_2 CB@1_mAd155_1 CB@1_mAd155_2 CB@1_mAd156_1 CB@1_mAd156_2 CB@1_mAd157_1 CB@1_mAd157_2 CB@1_mAd160_1 CB@1_mAd160_2 CB@1_mAd161_1 CB@1_mAd161_2 CB@1_mAd162_1 CB@1_mAd162_2 CB@1_mAd163_1 CB@1_mAd163_2 CB@1_mAd164_1 CB@1_mAd164_2 CB@1_mAd165_1 CB@1_mAd165_2 CB@1_mAd166_1 CB@1_mAd166_2 CB@1_mAd167_1 CB@1_mAd167_2 CB@1_mAd170_1 CB@1_mAd170_2 CB@1_mAd171_1 CB@1_mAd171_2 CB@1_mAd172_1 
+CB@1_mAd172_2 CB@1_mAd173_1 CB@1_mAd173_2 CB@1_mAd175_1 CB@1_mAd175_2 CB@1_mAd176_1 CB@1_mAd176_2 CB@1_mAd177_1 CB@1_mAd177_2 CB@1_mAd200_1 CB@1_mAd200_2 CB@1_mAd201_1 CB@1_mAd201_2 CB@1_mAd202_1 CB@1_mAd202_2 CB@1_mAd204_1 CB@1_mAd204_2 CB@1_mAd205_1 CB@1_mAd205_2 CB@1_mAd206_1 CB@1_mAd206_2 CB@1_mAd207_1 CB@1_mAd207_2 CB@1_mAd210_1 CB@1_mAd210_2 CB@1_mAd211_1 CB@1_mAd211_2 CB@1_mAd212_1 CB@1_mAd212_2 CB@1_mAd213_1 CB@1_mAd213_2 CB@1_mAd214_1 CB@1_mAd214_2 CB@1_mAd215_1 CB@1_mAd215_2 CB@1_mAd216_1 
+CB@1_mAd216_2 CB@1_mAd217_1 CB@1_mAd217_2 CB@1_mAd220_1 CB@1_mAd220_2 CB@1_mAd221_1 CB@1_mAd221_2 CB@1_mAd222_1 CB@1_mAd222_2 CB@1_mAd223_1 CB@1_mAd223_2 CB@1_mAd224_1 CB@1_mAd224_2 CB@1_mAd225_1 CB@1_mAd225_2 CB@1_mAd226_1 CB@1_mAd226_2 CB@1_mAd227_1 CB@1_mAd227_2 CB@1_mAd230_1 CB@1_mAd230_2 CB@1_mAd231_1 CB@1_mAd231_2 CB@1_mAd232_1 CB@1_mAd232_2 CB@1_mAd233_1 CB@1_mAd233_2 CB@1_mAd234_1 CB@1_mAd234_2 CB@1_mAd235_1 CB@1_mAd235_2 CB@1_mAd236_1 CB@1_mAd236_2 CB@1_mAd237_1 CB@1_mAd237_2 CB@1_mAd240_1 
+CB@1_mAd240_2 CB@1_mAd241_1 CB@1_mAd241_2 CB@1_mAd242_1 CB@1_mAd242_2 CB@1_mAd243_1 CB@1_mAd243_2 CB@1_mAd244_1 CB@1_mAd244_2 CB@1_mAd245_1 CB@1_mAd245_2 CB@1_mAd246_1 CB@1_mAd246_2 CB@1_mAd247_1 CB@1_mAd247_2 CB@1_mAd250_1 CB@1_mAd250_2 CB@1_mAd251_1 CB@1_mAd251_2 CB@1_mAd252_1 CB@1_mAd252_2 CB@1_mAd253_1 CB@1_mAd253_2 CB@1_mAd254_1 CB@1_mAd254_2 CB@1_mAd255_1 CB@1_mAd255_2 CB@1_mAd256_1 CB@1_mAd256_2 CB@1_mAd257_1 CB@1_mAd257_2 CB@1_mAd260_1 CB@1_mAd260_2 CB@1_mAd261_1 CB@1_mAd261_2 CB@1_mAd262_1 
+CB@1_mAd262_2 CB@1_mAd263_1 CB@1_mAd263_2 CB@1_mAd264_1 CB@1_mAd264_2 CB@1_mAd265_1 CB@1_mAd265_2 CB@1_mAd266_1 CB@1_mAd266_2 CB@1_mAd267_1 CB@1_mAd267_2 net@1459 net@1459 CB@1_mAd276_1 CB@1_mAd276_2 CB@1_mAd277_1 CB@1_mAd277_2 CB@1_mAd300_1 CB@1_mAd300_2 CB@1_mAd310_1 CB@1_mAd310_2 CB@1_mAd311_1 CB@1_mAd311_2 CB@1_mAd317_1 CB@1_mAd317_2 CB@1_mAd320_1 CB@1_mAd320_2 CB@1_mAd321_1 CB@1_mAd321_2 CB@1_mAd322_1 CB@1_mAd322_2 CB@1_mAd323_1 CB@1_mAd323_2 CB@1_mAd324_1 CB@1_mAd324_2 CB@1_mAd325_1 CB@1_mAd325_2 
+CB@1_mAd326_1 CB@1_mAd326_2 CB@1_mAd327_1 CB@1_mAd327_2 CB@1_mAd330_1 CB@1_mAd330_2 CB@1_mAd331_1 CB@1_mAd331_2 CB@1_mAd332_1 CB@1_mAd332_2 CB@1_mAd333_1 CB@1_mAd333_2 CB@1_mAd334_1 CB@1_mAd334_2 CB@1_mAd335_1 CB@1_mAd335_2 CB@1_mAd336_1 CB@1_mAd336_2 CB@1_mAd337_1 CB@1_mAd337_2 CB@1_mAd340_1 CB@1_mAd340_2 CB@1_mAd341_1 CB@1_mAd341_2 CB@1_mAd342_1 CB@1_mAd342_2 CB@1_mAd343_1 CB@1_mAd343_2 CB@1_mAd344_1 CB@1_mAd344_2 CB@1_mAd345_1 CB@1_mAd345_2 CB@1_mAd346_1 CB@1_mAd346_2 CB@1_mAd347_1 CB@1_mAd347_2 
+CB@1_mAd350_1 CB@1_mAd350_2 CB@1_mAd351_1 CB@1_mAd351_2 CB@1_mAd352_1 CB@1_mAd352_2 CB@1_mAd353_1 CB@1_mAd353_2 CB@1_mAd354_1 CB@1_mAd354_2 CB@1_mAd355_1 CB@1_mAd355_2 CB@1_mAd356_1 CB@1_mAd356_2 CB@1_mAd357_1 CB@1_mAd357_2 CB@1_mAd360_1 CB@1_mAd360_2 CB@1_mAd361_1 CB@1_mAd361_2 CB@1_mAd362_1 CB@1_mAd362_2 CB@1_mAd363_1 CB@1_mAd363_2 net@1460 net@1460 CB@1_mAd365_1 CB@1_mAd365_2 CB@1_mAd366_1 CB@1_mAd366_2 CB@1_mAd367_1 CB@1_mAd367_2 CB@1_mAd371_1 CB@1_mAd371_2 CB@1_mAd372_1 CB@1_mAd372_2 CB@1_mAd373_1 
+CB@1_mAd373_2 CB@1_mAd374_1 CB@1_mAd374_2 CB@1_mAd375_1 CB@1_mAd375_2 CB@1_mAd376_1 CB@1_mAd376_2 CB@1_mAd377_1 CB@1_mAd377_2 CB@1_mAd400_1 CB@1_mAd400_2 CB@1_mAd401_1 CB@1_mAd401_2 CB@1_mAd402_1 CB@1_mAd402_2 CB@1_mAd403_1 CB@1_mAd403_2 CB@1_mAd404_1 CB@1_mAd404_2 CB@1_mAd405_1 CB@1_mAd405_2 CB@1_mAd406_1 CB@1_mAd406_2 CB@1_mAd407_1 CB@1_mAd407_2 CB@1_mAd410_1 CB@1_mAd410_2 CB@1_mAd411_1 CB@1_mAd411_2 CB@1_mAd412_1 CB@1_mAd412_2 CB@1_mAd413_1 CB@1_mAd413_2 CB@1_mAd414_1 CB@1_mAd414_2 CB@1_mAd415_1 
+CB@1_mAd415_2 CB@1_mAd416_1 CB@1_mAd416_2 CB@1_mAd417_1 CB@1_mAd417_2 CB@1_mAd420_1 CB@1_mAd420_2 CB@1_mAd421_1 CB@1_mAd421_2 CB@1_mAd422_1 CB@1_mAd422_2 CB@1_mAd423_1 CB@1_mAd423_2 CB@1_mAd424_1 CB@1_mAd424_2 CB@1_mAd425_1 CB@1_mAd425_2 CB@1_mAd426_1 CB@1_mAd426_2 CB@1_mAd427_1 CB@1_mAd427_2 CB@1_mAd430_1 CB@1_mAd430_2 CB@1_mAd431_1 CB@1_mAd431_2 CB@1_mAd432_1 CB@1_mAd432_2 CB@1_mAd433_1 CB@1_mAd433_2 CB@1_mAd434_1 CB@1_mAd434_2 CB@1_mAd435_1 CB@1_mAd435_2 CB@1_mAd436_1 CB@1_mAd436_2 CB@1_mAd437_1 
+CB@1_mAd437_2 CB@1_mAd440_1 CB@1_mAd440_2 CB@1_mAd441_1 CB@1_mAd441_2 CB@1_mAd442_1 CB@1_mAd442_2 CB@1_mAd443_1 CB@1_mAd443_2 CB@1_mAd444_1 CB@1_mAd444_2 CB@1_mAd445_1 CB@1_mAd445_2 CB@1_mAd446_1 CB@1_mAd446_2 CB@1_mAd447_1 CB@1_mAd447_2 CB@1_mAd450_1 CB@1_mAd450_2 CB@1_mAd451_1 CB@1_mAd451_2 CB@1_mAd452_1 CB@1_mAd452_2 CB@1_mAd453_1 CB@1_mAd453_2 CB@1_mAd454_1 CB@1_mAd454_2 CB@1_mAd455_1 CB@1_mAd455_2 CB@1_mAd456_1 CB@1_mAd456_2 CB@1_mAd457_1 CB@1_mAd457_2 CB@1_mAd460_1 CB@1_mAd460_2 CB@1_mAd466_1 
+CB@1_mAd466_2 CB@1_mAd467_1 CB@1_mAd467_2 CB@1_mAd500_1 CB@1_mAd500_2 CB@1_mAd501_1 CB@1_mAd501_2 CB@1_mAd502_1 CB@1_mAd502_2 CB@1_mAd508_1 CB@1_mAd508_2 CB@1_mAd509_1 CB@1_mAd509_2 CB@1_mAd512_1 CB@1_mAd512_2 CB@1_mAd513_1 CB@1_mAd513_2 CB@1_mAd514_1 CB@1_mAd514_2 CB@1_mAd515_1 CB@1_mAd515_2 CB@1_mAd516_1 CB@1_mAd516_2 CB@1_mAd517_1 CB@1_mAd517_2 CB@1_mAd520_1 CB@1_mAd520_2 CB@1_mAd521_1 CB@1_mAd521_2 CB@1_mAd522_1 CB@1_mAd522_2 CB@1_mAd523_1 CB@1_mAd523_2 CB@1_mAd524_1 CB@1_mAd524_2 CB@1_mAd525_1 
+CB@1_mAd525_2 CB@1_mAd526_1 CB@1_mAd526_2 CB@1_mAd527_1 CB@1_mAd527_2 CB@1_mAd530_1 CB@1_mAd530_2 CB@1_mAd531_1 CB@1_mAd531_2 CB@1_mAd532_1 CB@1_mAd532_2 CB@1_mAd533_1 CB@1_mAd533_2 CB@1_mAd534_1 CB@1_mAd534_2 CB@1_mAd535_1 CB@1_mAd535_2 CB@1_mAd536_1 CB@1_mAd536_2 CB@1_mAd537_1 CB@1_mAd537_2 CB@1_mAd540_1 CB@1_mAd540_2 CB@1_mAd541_1 CB@1_mAd541_2 CB@1_mAd542_1 CB@1_mAd542_2 CB@1_mAd543_1 CB@1_mAd543_2 CB@1_mAd544_1 CB@1_mAd544_2 CB@1_mAd545_1 CB@1_mAd545_2 CB@1_mAd546_1 CB@1_mAd546_2 CB@1_mAd547_1 
+CB@1_mAd547_2 CB@1_mAd550_1 CB@1_mAd550_2 CB@1_mAd551_1 CB@1_mAd551_2 CB@1_mAd552_1 CB@1_mAd552_2 CB@1_mAd553_1 CB@1_mAd553_2 CB@1_mAd554_1 CB@1_mAd554_2 CB@1_mAd555_1 CB@1_mAd555_2 CB@1_mAd556_1 CB@1_mAd556_2 CB@1_mAd557_1 CB@1_mAd557_2 CB@1_mAd560_1 CB@1_mAd560_2 CB@1_mAd561_1 CB@1_mAd561_2 CB@1_mAd562_1 CB@1_mAd562_2 CB@1_mAd563_1 CB@1_mAd563_2 CB@1_mAd564_1 CB@1_mAd564_2 CB@1_mAd565_1 CB@1_mAd565_2 CB@1_mAd566_1 CB@1_mAd566_2 CB@1_mAd567_1 CB@1_mAd567_2 CB@1_mAd570_1 CB@1_mAd570_2 CB@1_mAd571_1 
+CB@1_mAd571_2 CB@1_mAd572_1 CB@1_mAd572_2 CB@1_mAd573_1 CB@1_mAd573_2 CB@1_mAd575_1 CB@1_mAd575_2 CB@1_mAd576_1 CB@1_mAd576_2 CB@1_mAd577_1 CB@1_mAd577_2 CB@1_mAd600_1 CB@1_mAd600_2 CB@1_mAd601_1 CB@1_mAd601_2 CB@1_mAd602_1 CB@1_mAd602_2 CB@1_mAd604_1 CB@1_mAd604_2 CB@1_mAd605_1 CB@1_mAd605_2 CB@1_mAd606_1 CB@1_mAd606_2 CB@1_mAd607_1 CB@1_mAd607_2 CB@1_mAd610_1 CB@1_mAd610_2 CB@1_mAd611_1 CB@1_mAd611_2 CB@1_mAd612_1 CB@1_mAd612_2 CB@1_mAd613_1 CB@1_mAd613_2 CB@1_mAd614_1 CB@1_mAd614_2 CB@1_mAd615_1 
+CB@1_mAd615_2 CB@1_mAd616_1 CB@1_mAd616_2 CB@1_mAd617_1 CB@1_mAd617_2 CB@1_mAd620_1 CB@1_mAd620_2 CB@1_mAd621_1 CB@1_mAd621_2 CB@1_mAd622_1 CB@1_mAd622_2 CB@1_mAd623_1 CB@1_mAd623_2 CB@1_mAd624_1 CB@1_mAd624_2 CB@1_mAd625_1 CB@1_mAd625_2 CB@1_mAd626_1 CB@1_mAd626_2 CB@1_mAd627_1 CB@1_mAd627_2 CB@1_mAd630_1 CB@1_mAd630_2 CB@1_mAd631_1 CB@1_mAd631_2 CB@1_mAd632_1 CB@1_mAd632_2 CB@1_mAd633_1 CB@1_mAd633_2 CB@1_mAd634_1 CB@1_mAd634_2 CB@1_mAd635_1 CB@1_mAd635_2 CB@1_mAd636_1 CB@1_mAd636_2 CB@1_mAd637_1 
+CB@1_mAd637_2 CB@1_mAd640_1 CB@1_mAd640_2 CB@1_mAd641_1 CB@1_mAd641_2 CB@1_mAd642_1 CB@1_mAd642_2 CB@1_mAd643_1 CB@1_mAd643_2 CB@1_mAd644_1 CB@1_mAd644_2 CB@1_mAd645_1 CB@1_mAd645_2 CB@1_mAd646_1 CB@1_mAd646_2 CB@1_mAd647_1 CB@1_mAd647_2 CB@1_mAd650_1 CB@1_mAd650_2 CB@1_mAd651_1 CB@1_mAd651_2 CB@1_mAd652_1 CB@1_mAd652_2 CB@1_mAd653_1 CB@1_mAd653_2 CB@1_mAd654_1 CB@1_mAd654_2 CB@1_mAd655_1 CB@1_mAd655_2 CB@1_mAd656_1 CB@1_mAd656_2 CB@1_mAd657_1 CB@1_mAd657_2 CB@1_mAd660_1 CB@1_mAd660_2 CB@1_mAd661_1 
+CB@1_mAd661_2 CB@1_mAd662_1 CB@1_mAd662_2 CB@1_mAd663_1 CB@1_mAd663_2 CB@1_mAd664_1 CB@1_mAd664_2 CB@1_mAd665_1 CB@1_mAd665_2 CB@1_mAd666_1 CB@1_mAd666_2 CB@1_mAd667_1 CB@1_mAd667_2 CB@1_mAd675_1 CB@1_mAd675_2 CB@1_mAd676_1 CB@1_mAd676_2 CB@1_mAd677_1 CB@1_mAd677_2 CB@1_mAd700_1 CB@1_mAd700_2 CB@1_mAd710_1 CB@1_mAd710_2 CB@1_mAd711_1 CB@1_mAd711_2 CB@1_mAd717_1 CB@1_mAd717_2 CB@1_mAd720_1 CB@1_mAd720_2 CB@1_mAd721_1 CB@1_mAd721_2 CB@1_mAd722_1 CB@1_mAd722_2 CB@1_mAd723_1 CB@1_mAd723_2 CB@1_mAd724_1 
+CB@1_mAd724_2 CB@1_mAd725_1 CB@1_mAd725_2 CB@1_mAd726_1 CB@1_mAd726_2 CB@1_mAd727_1 CB@1_mAd727_2 CB@1_mAd730_1 CB@1_mAd730_2 CB@1_mAd731_1 CB@1_mAd731_2 CB@1_mAd732_1 CB@1_mAd732_2 CB@1_mAd733_1 CB@1_mAd733_2 CB@1_mAd734_1 CB@1_mAd734_2 CB@1_mAd735_1 CB@1_mAd735_2 CB@1_mAd736_1 CB@1_mAd736_2 CB@1_mAd737_1 CB@1_mAd737_2 CB@1_mAd740_1 CB@1_mAd740_2 CB@1_mAd741_1 CB@1_mAd741_2 CB@1_mAd742_1 CB@1_mAd742_2 CB@1_mAd743_1 CB@1_mAd743_2 CB@1_mAd744_1 CB@1_mAd744_2 CB@1_mAd745_1 CB@1_mAd745_2 CB@1_mAd746_1 
+CB@1_mAd746_2 CB@1_mAd747_1 CB@1_mAd747_2 CB@1_mAd750_1 CB@1_mAd750_2 CB@1_mAd751_1 CB@1_mAd751_2 CB@1_mAd752_1 CB@1_mAd752_2 CB@1_mAd753_1 CB@1_mAd753_2 CB@1_mAd754_1 CB@1_mAd754_2 CB@1_mAd755_1 CB@1_mAd755_2 CB@1_mAd756_1 CB@1_mAd756_2 CB@1_mAd757_1 CB@1_mAd757_2 CB@1_mAd760_1 CB@1_mAd760_2 CB@1_mAd761_1 CB@1_mAd761_2 CB@1_mAd762_1 CB@1_mAd762_2 CB@1_mAd763_1 CB@1_mAd763_2 CB@1_mAd764_1 CB@1_mAd764_2 CB@1_mAd765_1 CB@1_mAd765_2 CB@1_mAd766_1 CB@1_mAd766_2 CB@1_mAd767_1 CB@1_mAd767_2 CB@1_mAd771_1 
+CB@1_mAd771_2 CB@1_mAd772_1 CB@1_mAd772_2 CB@1_mAd773_1 CB@1_mAd773_2 CB@1_mAd774_1 CB@1_mAd774_2 CB@1_mAd775_1 CB@1_mAd775_2 CB@1_mAd776_1 CB@1_mAd776_2 CB@1_mAd777_1 CB@1_mAd777_2 CB@1_X0 CB@1_X1 CB@1_X10 CB@1_X11 CB@1_X12 CB@1_X13 CB@1_X2 net@1447 CB@1_X4 CB@1_X5 CB@1_X6 CB@1_X7 CB@1_X8 CB@1_X9 CB@1_Y1 CB@1_Y10 CB@1_Y11 CB@1_Y12 CB@1_Y2 CB@1_Y3 CB@1_Y4 CB@1_Y5 CB@1_Y6 CB@1_Y7 CB@1_Y8 CB@1_Y9 CB@1_Z1 CB@1_Z10 CB@1_Z11 CB@1_Z12 out2 out1 CB@1_Z4 CB@1_Z5 CB@1_Z6 CB@1_Z7 CB@1_Z8 CB@1_Z9 _5400TP094__CB
XCB@2 CB@2_K0 CB@2_K1 CB@2_K10 CB@2_K11 CB@2_K12 CB@2_K13 CB@2_K2 CB@2_K3 CB@2_K4 CB@2_K5 CB@2_K6 CB@2_K7 CB@2_K8 CB@2_K9 CB@2_mAd000_1 CB@2_mAd000_2 CB@2_mAd001_1 CB@2_mAd001_2 CB@2_mAd002_1 CB@2_mAd002_2 CB@2_mAd003_1 CB@2_mAd003_2 CB@2_mAd004_1 CB@2_mAd004_2 CB@2_mAd005_1 CB@2_mAd005_2 CB@2_mAd006_1 CB@2_mAd006_2 CB@2_mAd007_1 CB@2_mAd007_2 CB@2_mAd010_1 CB@2_mAd010_2 CB@2_mAd011_1 CB@2_mAd011_2 CB@2_mAd012_1 CB@2_mAd012_2 CB@2_mAd013_1 CB@2_mAd013_2 CB@2_mAd014_1 CB@2_mAd014_2 CB@2_mAd015_1 
+CB@2_mAd015_2 CB@2_mAd016_1 CB@2_mAd016_2 CB@2_mAd017_1 CB@2_mAd017_2 CB@2_mAd020_1 CB@2_mAd020_2 CB@2_mAd021_1 CB@2_mAd021_2 CB@2_mAd022_1 CB@2_mAd022_2 CB@2_mAd023_1 CB@2_mAd023_2 CB@2_mAd024_1 CB@2_mAd024_2 CB@2_mAd025_1 CB@2_mAd025_2 CB@2_mAd026_1 CB@2_mAd026_2 CB@2_mAd027_1 CB@2_mAd027_2 CB@2_mAd030_1 CB@2_mAd030_2 CB@2_mAd031_1 CB@2_mAd031_2 CB@2_mAd032_1 CB@2_mAd032_2 CB@2_mAd033_1 CB@2_mAd033_2 CB@2_mAd034_1 CB@2_mAd034_2 CB@2_mAd035_1 CB@2_mAd035_2 CB@2_mAd036_1 CB@2_mAd036_2 CB@2_mAd037_1 
+CB@2_mAd037_2 CB@2_mAd040_1 CB@2_mAd040_2 CB@2_mAd041_1 CB@2_mAd041_2 CB@2_mAd042_1 CB@2_mAd042_2 CB@2_mAd043_1 CB@2_mAd043_2 CB@2_mAd044_1 CB@2_mAd044_2 CB@2_mAd045_1 CB@2_mAd045_2 CB@2_mAd046_1 CB@2_mAd046_2 CB@2_mAd047_1 CB@2_mAd047_2 CB@2_mAd050_1 CB@2_mAd050_2 CB@2_mAd051_1 CB@2_mAd051_2 CB@2_mAd052_1 CB@2_mAd052_2 CB@2_mAd053_1 CB@2_mAd053_2 CB@2_mAd054_1 CB@2_mAd054_2 CB@2_mAd055_1 CB@2_mAd055_2 CB@2_mAd056_1 CB@2_mAd056_2 CB@2_mAd057_1 CB@2_mAd057_2 CB@2_mAd060_1 CB@2_mAd060_2 CB@2_mAd066_1 
+CB@2_mAd066_2 CB@2_mAd067_1 CB@2_mAd067_2 CB@2_mAd100_1 CB@2_mAd100_2 CB@2_mAd101_1 CB@2_mAd101_2 CB@2_mAd102_1 CB@2_mAd102_2 CB@2_mAd110_1 CB@2_mAd110_2 CB@2_mAd111_1 CB@2_mAd111_2 CB@2_mAd112_1 CB@2_mAd112_2 CB@2_mAd113_1 CB@2_mAd113_2 CB@2_mAd114_1 CB@2_mAd114_2 CB@2_mAd115_1 CB@2_mAd115_2 CB@2_mAd116_1 CB@2_mAd116_2 CB@2_mAd117_1 CB@2_mAd117_2 CB@2_mAd120_1 CB@2_mAd120_2 CB@2_mAd121_1 CB@2_mAd121_2 CB@2_mAd122_1 CB@2_mAd122_2 CB@2_mAd123_1 CB@2_mAd123_2 CB@2_mAd124_1 CB@2_mAd124_2 CB@2_mAd125_1 
+CB@2_mAd125_2 CB@2_mAd126_1 CB@2_mAd126_2 CB@2_mAd127_1 CB@2_mAd127_2 CB@2_mAd130_1 CB@2_mAd130_2 CB@2_mAd131_1 CB@2_mAd131_2 CB@2_mAd132_1 CB@2_mAd132_2 CB@2_mAd133_1 CB@2_mAd133_2 CB@2_mAd134_1 CB@2_mAd134_2 CB@2_mAd135_1 CB@2_mAd135_2 CB@2_mAd136_1 CB@2_mAd136_2 CB@2_mAd137_1 CB@2_mAd137_2 CB@2_mAd140_1 CB@2_mAd140_2 CB@2_mAd141_1 CB@2_mAd141_2 CB@2_mAd142_1 CB@2_mAd142_2 CB@2_mAd143_1 CB@2_mAd143_2 CB@2_mAd144_1 CB@2_mAd144_2 CB@2_mAd145_1 CB@2_mAd145_2 CB@2_mAd146_1 CB@2_mAd146_2 CB@2_mAd147_1 
+CB@2_mAd147_2 CB@2_mAd150_1 CB@2_mAd150_2 CB@2_mAd151_1 CB@2_mAd151_2 CB@2_mAd152_1 CB@2_mAd152_2 CB@2_mAd153_1 CB@2_mAd153_2 CB@2_mAd154_1 CB@2_mAd154_2 CB@2_mAd155_1 CB@2_mAd155_2 CB@2_mAd156_1 CB@2_mAd156_2 CB@2_mAd157_1 CB@2_mAd157_2 CB@2_mAd160_1 CB@2_mAd160_2 CB@2_mAd161_1 CB@2_mAd161_2 CB@2_mAd162_1 CB@2_mAd162_2 CB@2_mAd163_1 CB@2_mAd163_2 CB@2_mAd164_1 CB@2_mAd164_2 CB@2_mAd165_1 CB@2_mAd165_2 CB@2_mAd166_1 CB@2_mAd166_2 CB@2_mAd167_1 CB@2_mAd167_2 CB@2_mAd170_1 CB@2_mAd170_2 CB@2_mAd171_1 
+CB@2_mAd171_2 CB@2_mAd172_1 CB@2_mAd172_2 CB@2_mAd173_1 CB@2_mAd173_2 CB@2_mAd175_1 CB@2_mAd175_2 CB@2_mAd176_1 CB@2_mAd176_2 CB@2_mAd177_1 CB@2_mAd177_2 CB@2_mAd200_1 CB@2_mAd200_2 CB@2_mAd201_1 CB@2_mAd201_2 CB@2_mAd202_1 CB@2_mAd202_2 CB@2_mAd204_1 CB@2_mAd204_2 CB@2_mAd205_1 CB@2_mAd205_2 CB@2_mAd206_1 CB@2_mAd206_2 CB@2_mAd207_1 CB@2_mAd207_2 CB@2_mAd210_1 CB@2_mAd210_2 CB@2_mAd211_1 CB@2_mAd211_2 CB@2_mAd212_1 CB@2_mAd212_2 CB@2_mAd213_1 CB@2_mAd213_2 CB@2_mAd214_1 CB@2_mAd214_2 CB@2_mAd215_1 
+CB@2_mAd215_2 CB@2_mAd216_1 CB@2_mAd216_2 CB@2_mAd217_1 CB@2_mAd217_2 CB@2_mAd220_1 CB@2_mAd220_2 CB@2_mAd221_1 CB@2_mAd221_2 CB@2_mAd222_1 CB@2_mAd222_2 CB@2_mAd223_1 CB@2_mAd223_2 CB@2_mAd224_1 CB@2_mAd224_2 CB@2_mAd225_1 CB@2_mAd225_2 CB@2_mAd226_1 CB@2_mAd226_2 CB@2_mAd227_1 CB@2_mAd227_2 CB@2_mAd230_1 CB@2_mAd230_2 CB@2_mAd231_1 CB@2_mAd231_2 CB@2_mAd232_1 CB@2_mAd232_2 CB@2_mAd233_1 CB@2_mAd233_2 CB@2_mAd234_1 CB@2_mAd234_2 CB@2_mAd235_1 CB@2_mAd235_2 CB@2_mAd236_1 CB@2_mAd236_2 CB@2_mAd237_1 
+CB@2_mAd237_2 CB@2_mAd240_1 CB@2_mAd240_2 CB@2_mAd241_1 CB@2_mAd241_2 CB@2_mAd242_1 CB@2_mAd242_2 CB@2_mAd243_1 CB@2_mAd243_2 CB@2_mAd244_1 CB@2_mAd244_2 CB@2_mAd245_1 CB@2_mAd245_2 CB@2_mAd246_1 CB@2_mAd246_2 CB@2_mAd247_1 CB@2_mAd247_2 CB@2_mAd250_1 CB@2_mAd250_2 CB@2_mAd251_1 CB@2_mAd251_2 CB@2_mAd252_1 CB@2_mAd252_2 CB@2_mAd253_1 CB@2_mAd253_2 CB@2_mAd254_1 CB@2_mAd254_2 CB@2_mAd255_1 CB@2_mAd255_2 CB@2_mAd256_1 CB@2_mAd256_2 CB@2_mAd257_1 CB@2_mAd257_2 CB@2_mAd260_1 CB@2_mAd260_2 CB@2_mAd261_1 
+CB@2_mAd261_2 CB@2_mAd262_1 CB@2_mAd262_2 CB@2_mAd263_1 CB@2_mAd263_2 CB@2_mAd264_1 CB@2_mAd264_2 CB@2_mAd265_1 CB@2_mAd265_2 CB@2_mAd266_1 CB@2_mAd266_2 CB@2_mAd267_1 CB@2_mAd267_2 CB@2_mAd275_1 CB@2_mAd275_2 CB@2_mAd276_1 CB@2_mAd276_2 CB@2_mAd277_1 CB@2_mAd277_2 CB@2_mAd300_1 CB@2_mAd300_2 CB@2_mAd310_1 CB@2_mAd310_2 CB@2_mAd311_1 CB@2_mAd311_2 CB@2_mAd317_1 CB@2_mAd317_2 CB@2_mAd320_1 CB@2_mAd320_2 CB@2_mAd321_1 CB@2_mAd321_2 CB@2_mAd322_1 CB@2_mAd322_2 CB@2_mAd323_1 CB@2_mAd323_2 CB@2_mAd324_1 
+CB@2_mAd324_2 CB@2_mAd325_1 CB@2_mAd325_2 CB@2_mAd326_1 CB@2_mAd326_2 CB@2_mAd327_1 CB@2_mAd327_2 CB@2_mAd330_1 CB@2_mAd330_2 CB@2_mAd331_1 CB@2_mAd331_2 CB@2_mAd332_1 CB@2_mAd332_2 CB@2_mAd333_1 CB@2_mAd333_2 CB@2_mAd334_1 CB@2_mAd334_2 CB@2_mAd335_1 CB@2_mAd335_2 CB@2_mAd336_1 CB@2_mAd336_2 CB@2_mAd337_1 CB@2_mAd337_2 CB@2_mAd340_1 CB@2_mAd340_2 CB@2_mAd341_1 CB@2_mAd341_2 CB@2_mAd342_1 CB@2_mAd342_2 CB@2_mAd343_1 CB@2_mAd343_2 CB@2_mAd344_1 CB@2_mAd344_2 CB@2_mAd345_1 CB@2_mAd345_2 CB@2_mAd346_1 
+CB@2_mAd346_2 CB@2_mAd347_1 CB@2_mAd347_2 CB@2_mAd350_1 CB@2_mAd350_2 CB@2_mAd351_1 CB@2_mAd351_2 CB@2_mAd352_1 CB@2_mAd352_2 CB@2_mAd353_1 CB@2_mAd353_2 CB@2_mAd354_1 CB@2_mAd354_2 CB@2_mAd355_1 CB@2_mAd355_2 CB@2_mAd356_1 CB@2_mAd356_2 CB@2_mAd357_1 CB@2_mAd357_2 CB@2_mAd360_1 CB@2_mAd360_2 CB@2_mAd361_1 CB@2_mAd361_2 CB@2_mAd362_1 CB@2_mAd362_2 CB@2_mAd363_1 CB@2_mAd363_2 CB@2_mAd364_1 CB@2_mAd364_2 CB@2_mAd365_1 CB@2_mAd365_2 CB@2_mAd366_1 CB@2_mAd366_2 CB@2_mAd367_1 CB@2_mAd367_2 CB@2_mAd371_1 
+CB@2_mAd371_2 CB@2_mAd372_1 CB@2_mAd372_2 CB@2_mAd373_1 CB@2_mAd373_2 CB@2_mAd374_1 CB@2_mAd374_2 CB@2_mAd375_1 CB@2_mAd375_2 CB@2_mAd376_1 CB@2_mAd376_2 CB@2_mAd377_1 CB@2_mAd377_2 CB@2_mAd400_1 CB@2_mAd400_2 CB@2_mAd401_1 CB@2_mAd401_2 CB@2_mAd402_1 CB@2_mAd402_2 CB@2_mAd403_1 CB@2_mAd403_2 CB@2_mAd404_1 CB@2_mAd404_2 CB@2_mAd405_1 CB@2_mAd405_2 CB@2_mAd406_1 CB@2_mAd406_2 CB@2_mAd407_1 CB@2_mAd407_2 CB@2_mAd410_1 CB@2_mAd410_2 CB@2_mAd411_1 CB@2_mAd411_2 CB@2_mAd412_1 CB@2_mAd412_2 CB@2_mAd413_1 
+CB@2_mAd413_2 CB@2_mAd414_1 CB@2_mAd414_2 CB@2_mAd415_1 CB@2_mAd415_2 CB@2_mAd416_1 CB@2_mAd416_2 CB@2_mAd417_1 CB@2_mAd417_2 CB@2_mAd420_1 CB@2_mAd420_2 CB@2_mAd421_1 CB@2_mAd421_2 CB@2_mAd422_1 CB@2_mAd422_2 CB@2_mAd423_1 CB@2_mAd423_2 CB@2_mAd424_1 CB@2_mAd424_2 CB@2_mAd425_1 CB@2_mAd425_2 CB@2_mAd426_1 CB@2_mAd426_2 CB@2_mAd427_1 CB@2_mAd427_2 CB@2_mAd430_1 CB@2_mAd430_2 CB@2_mAd431_1 CB@2_mAd431_2 CB@2_mAd432_1 CB@2_mAd432_2 CB@2_mAd433_1 CB@2_mAd433_2 CB@2_mAd434_1 CB@2_mAd434_2 CB@2_mAd435_1 
+CB@2_mAd435_2 CB@2_mAd436_1 CB@2_mAd436_2 CB@2_mAd437_1 CB@2_mAd437_2 CB@2_mAd440_1 CB@2_mAd440_2 CB@2_mAd441_1 CB@2_mAd441_2 CB@2_mAd442_1 CB@2_mAd442_2 CB@2_mAd443_1 CB@2_mAd443_2 CB@2_mAd444_1 CB@2_mAd444_2 CB@2_mAd445_1 CB@2_mAd445_2 CB@2_mAd446_1 CB@2_mAd446_2 CB@2_mAd447_1 CB@2_mAd447_2 CB@2_mAd450_1 CB@2_mAd450_2 CB@2_mAd451_1 CB@2_mAd451_2 CB@2_mAd452_1 CB@2_mAd452_2 CB@2_mAd453_1 CB@2_mAd453_2 CB@2_mAd454_1 CB@2_mAd454_2 CB@2_mAd455_1 CB@2_mAd455_2 CB@2_mAd456_1 CB@2_mAd456_2 CB@2_mAd457_1 
+CB@2_mAd457_2 CB@2_mAd460_1 CB@2_mAd460_2 CB@2_mAd466_1 CB@2_mAd466_2 CB@2_mAd467_1 CB@2_mAd467_2 CB@2_mAd500_1 CB@2_mAd500_2 CB@2_mAd501_1 CB@2_mAd501_2 CB@2_mAd502_1 CB@2_mAd502_2 CB@2_mAd508_1 CB@2_mAd508_2 CB@2_mAd509_1 CB@2_mAd509_2 CB@2_mAd512_1 CB@2_mAd512_2 CB@2_mAd513_1 CB@2_mAd513_2 CB@2_mAd514_1 CB@2_mAd514_2 CB@2_mAd515_1 CB@2_mAd515_2 CB@2_mAd516_1 CB@2_mAd516_2 CB@2_mAd517_1 CB@2_mAd517_2 CB@2_mAd520_1 CB@2_mAd520_2 CB@2_mAd521_1 CB@2_mAd521_2 CB@2_mAd522_1 CB@2_mAd522_2 CB@2_mAd523_1 
+CB@2_mAd523_2 CB@2_mAd524_1 CB@2_mAd524_2 CB@2_mAd525_1 CB@2_mAd525_2 CB@2_mAd526_1 CB@2_mAd526_2 CB@2_mAd527_1 CB@2_mAd527_2 CB@2_mAd530_1 CB@2_mAd530_2 CB@2_mAd531_1 CB@2_mAd531_2 CB@2_mAd532_1 CB@2_mAd532_2 CB@2_mAd533_1 CB@2_mAd533_2 CB@2_mAd534_1 CB@2_mAd534_2 CB@2_mAd535_1 CB@2_mAd535_2 CB@2_mAd536_1 CB@2_mAd536_2 CB@2_mAd537_1 CB@2_mAd537_2 CB@2_mAd540_1 CB@2_mAd540_2 CB@2_mAd541_1 CB@2_mAd541_2 CB@2_mAd542_1 CB@2_mAd542_2 CB@2_mAd543_1 CB@2_mAd543_2 CB@2_mAd544_1 CB@2_mAd544_2 CB@2_mAd545_1 
+CB@2_mAd545_2 CB@2_mAd546_1 CB@2_mAd546_2 CB@2_mAd547_1 CB@2_mAd547_2 CB@2_mAd550_1 CB@2_mAd550_2 CB@2_mAd551_1 CB@2_mAd551_2 CB@2_mAd552_1 CB@2_mAd552_2 CB@2_mAd553_1 CB@2_mAd553_2 CB@2_mAd554_1 CB@2_mAd554_2 CB@2_mAd555_1 CB@2_mAd555_2 CB@2_mAd556_1 CB@2_mAd556_2 CB@2_mAd557_1 CB@2_mAd557_2 CB@2_mAd560_1 CB@2_mAd560_2 CB@2_mAd561_1 CB@2_mAd561_2 CB@2_mAd562_1 CB@2_mAd562_2 CB@2_mAd563_1 CB@2_mAd563_2 CB@2_mAd564_1 CB@2_mAd564_2 CB@2_mAd565_1 CB@2_mAd565_2 CB@2_mAd566_1 CB@2_mAd566_2 CB@2_mAd567_1 
+CB@2_mAd567_2 CB@2_mAd570_1 CB@2_mAd570_2 CB@2_mAd571_1 CB@2_mAd571_2 CB@2_mAd572_1 CB@2_mAd572_2 CB@2_mAd573_1 CB@2_mAd573_2 CB@2_mAd575_1 CB@2_mAd575_2 CB@2_mAd576_1 CB@2_mAd576_2 CB@2_mAd577_1 CB@2_mAd577_2 CB@2_mAd600_1 CB@2_mAd600_2 CB@2_mAd601_1 CB@2_mAd601_2 CB@2_mAd602_1 CB@2_mAd602_2 CB@2_mAd604_1 CB@2_mAd604_2 CB@2_mAd605_1 CB@2_mAd605_2 CB@2_mAd606_1 CB@2_mAd606_2 CB@2_mAd607_1 CB@2_mAd607_2 CB@2_mAd610_1 CB@2_mAd610_2 CB@2_mAd611_1 CB@2_mAd611_2 CB@2_mAd612_1 CB@2_mAd612_2 CB@2_mAd613_1 
+CB@2_mAd613_2 CB@2_mAd614_1 CB@2_mAd614_2 CB@2_mAd615_1 CB@2_mAd615_2 CB@2_mAd616_1 CB@2_mAd616_2 CB@2_mAd617_1 CB@2_mAd617_2 CB@2_mAd620_1 CB@2_mAd620_2 CB@2_mAd621_1 CB@2_mAd621_2 CB@2_mAd622_1 CB@2_mAd622_2 CB@2_mAd623_1 CB@2_mAd623_2 CB@2_mAd624_1 CB@2_mAd624_2 CB@2_mAd625_1 CB@2_mAd625_2 CB@2_mAd626_1 CB@2_mAd626_2 CB@2_mAd627_1 CB@2_mAd627_2 CB@2_mAd630_1 CB@2_mAd630_2 CB@2_mAd631_1 CB@2_mAd631_2 CB@2_mAd632_1 CB@2_mAd632_2 CB@2_mAd633_1 CB@2_mAd633_2 CB@2_mAd634_1 CB@2_mAd634_2 CB@2_mAd635_1 
+CB@2_mAd635_2 CB@2_mAd636_1 CB@2_mAd636_2 CB@2_mAd637_1 CB@2_mAd637_2 CB@2_mAd640_1 CB@2_mAd640_2 CB@2_mAd641_1 CB@2_mAd641_2 CB@2_mAd642_1 CB@2_mAd642_2 CB@2_mAd643_1 CB@2_mAd643_2 CB@2_mAd644_1 CB@2_mAd644_2 CB@2_mAd645_1 CB@2_mAd645_2 CB@2_mAd646_1 CB@2_mAd646_2 CB@2_mAd647_1 CB@2_mAd647_2 CB@2_mAd650_1 CB@2_mAd650_2 CB@2_mAd651_1 CB@2_mAd651_2 CB@2_mAd652_1 CB@2_mAd652_2 CB@2_mAd653_1 CB@2_mAd653_2 CB@2_mAd654_1 CB@2_mAd654_2 CB@2_mAd655_1 CB@2_mAd655_2 CB@2_mAd656_1 CB@2_mAd656_2 CB@2_mAd657_1 
+CB@2_mAd657_2 CB@2_mAd660_1 CB@2_mAd660_2 CB@2_mAd661_1 CB@2_mAd661_2 CB@2_mAd662_1 CB@2_mAd662_2 CB@2_mAd663_1 CB@2_mAd663_2 CB@2_mAd664_1 CB@2_mAd664_2 CB@2_mAd665_1 CB@2_mAd665_2 CB@2_mAd666_1 CB@2_mAd666_2 CB@2_mAd667_1 CB@2_mAd667_2 CB@2_mAd675_1 CB@2_mAd675_2 CB@2_mAd676_1 CB@2_mAd676_2 CB@2_mAd677_1 CB@2_mAd677_2 CB@2_mAd700_1 CB@2_mAd700_2 CB@2_mAd710_1 CB@2_mAd710_2 CB@2_mAd711_1 CB@2_mAd711_2 CB@2_mAd717_1 CB@2_mAd717_2 CB@2_mAd720_1 CB@2_mAd720_2 CB@2_mAd721_1 CB@2_mAd721_2 CB@2_mAd722_1 
+CB@2_mAd722_2 CB@2_mAd723_1 CB@2_mAd723_2 CB@2_mAd724_1 CB@2_mAd724_2 CB@2_mAd725_1 CB@2_mAd725_2 CB@2_mAd726_1 CB@2_mAd726_2 CB@2_mAd727_1 CB@2_mAd727_2 CB@2_mAd730_1 CB@2_mAd730_2 CB@2_mAd731_1 CB@2_mAd731_2 CB@2_mAd732_1 CB@2_mAd732_2 CB@2_mAd733_1 CB@2_mAd733_2 CB@2_mAd734_1 CB@2_mAd734_2 CB@2_mAd735_1 CB@2_mAd735_2 CB@2_mAd736_1 CB@2_mAd736_2 CB@2_mAd737_1 CB@2_mAd737_2 CB@2_mAd740_1 CB@2_mAd740_2 CB@2_mAd741_1 CB@2_mAd741_2 CB@2_mAd742_1 CB@2_mAd742_2 CB@2_mAd743_1 CB@2_mAd743_2 CB@2_mAd744_1 
+CB@2_mAd744_2 CB@2_mAd745_1 CB@2_mAd745_2 CB@2_mAd746_1 CB@2_mAd746_2 CB@2_mAd747_1 CB@2_mAd747_2 CB@2_mAd750_1 CB@2_mAd750_2 CB@2_mAd751_1 CB@2_mAd751_2 CB@2_mAd752_1 CB@2_mAd752_2 CB@2_mAd753_1 CB@2_mAd753_2 CB@2_mAd754_1 CB@2_mAd754_2 CB@2_mAd755_1 CB@2_mAd755_2 CB@2_mAd756_1 CB@2_mAd756_2 CB@2_mAd757_1 CB@2_mAd757_2 CB@2_mAd760_1 CB@2_mAd760_2 CB@2_mAd761_1 CB@2_mAd761_2 CB@2_mAd762_1 CB@2_mAd762_2 CB@2_mAd763_1 CB@2_mAd763_2 CB@2_mAd764_1 CB@2_mAd764_2 CB@2_mAd765_1 CB@2_mAd765_2 CB@2_mAd766_1 
+CB@2_mAd766_2 CB@2_mAd767_1 CB@2_mAd767_2 CB@2_mAd771_1 CB@2_mAd771_2 CB@2_mAd772_1 CB@2_mAd772_2 CB@2_mAd773_1 CB@2_mAd773_2 CB@2_mAd774_1 CB@2_mAd774_2 CB@2_mAd775_1 CB@2_mAd775_2 CB@2_mAd776_1 CB@2_mAd776_2 CB@2_mAd777_1 CB@2_mAd777_2 CB@2_X0 CB@2_X1 CB@2_X10 CB@2_X11 CB@2_X12 CB@2_X13 CB@2_X2 CB@2_X3 CB@2_X4 CB@2_X5 CB@2_X6 CB@2_X7 CB@2_X8 CB@2_X9 CB@2_Y1 CB@2_Y10 CB@2_Y11 CB@2_Y12 CB@2_Y2 CB@2_Y3 CB@2_Y4 CB@2_Y5 CB@2_Y6 CB@2_Y7 CB@2_Y8 CB@2_Y9 CB@2_Z1 CB@2_Z10 CB@2_Z11 CB@2_Z12 CB@2_Z2 CB@2_Z3 CB@2_Z4 
+CB@2_Z5 CB@2_Z6 CB@2_Z7 CB@2_Z8 CB@2_Z9 _5400TP094__CB
XCB@3 CB@3_K0 CB@3_K1 CB@3_K10 CB@3_K11 CB@3_K12 CB@3_K13 CB@3_K2 CB@3_K3 CB@3_K4 CB@3_K5 CB@3_K6 CB@3_K7 CB@3_K8 CB@3_K9 CB@3_mAd000_1 CB@3_mAd000_2 CB@3_mAd001_1 CB@3_mAd001_2 CB@3_mAd002_1 CB@3_mAd002_2 CB@3_mAd003_1 CB@3_mAd003_2 CB@3_mAd004_1 CB@3_mAd004_2 CB@3_mAd005_1 CB@3_mAd005_2 CB@3_mAd006_1 CB@3_mAd006_2 CB@3_mAd007_1 CB@3_mAd007_2 CB@3_mAd010_1 CB@3_mAd010_2 CB@3_mAd011_1 CB@3_mAd011_2 CB@3_mAd012_1 CB@3_mAd012_2 CB@3_mAd013_1 CB@3_mAd013_2 CB@3_mAd014_1 CB@3_mAd014_2 CB@3_mAd015_1 
+CB@3_mAd015_2 CB@3_mAd016_1 CB@3_mAd016_2 CB@3_mAd017_1 CB@3_mAd017_2 CB@3_mAd020_1 CB@3_mAd020_2 CB@3_mAd021_1 CB@3_mAd021_2 CB@3_mAd022_1 CB@3_mAd022_2 CB@3_mAd023_1 CB@3_mAd023_2 CB@3_mAd024_1 CB@3_mAd024_2 CB@3_mAd025_1 CB@3_mAd025_2 CB@3_mAd026_1 CB@3_mAd026_2 CB@3_mAd027_1 CB@3_mAd027_2 CB@3_mAd030_1 CB@3_mAd030_2 CB@3_mAd031_1 CB@3_mAd031_2 CB@3_mAd032_1 CB@3_mAd032_2 CB@3_mAd033_1 CB@3_mAd033_2 CB@3_mAd034_1 CB@3_mAd034_2 CB@3_mAd035_1 CB@3_mAd035_2 CB@3_mAd036_1 CB@3_mAd036_2 CB@3_mAd037_1 
+CB@3_mAd037_2 CB@3_mAd040_1 CB@3_mAd040_2 CB@3_mAd041_1 CB@3_mAd041_2 CB@3_mAd042_1 CB@3_mAd042_2 CB@3_mAd043_1 CB@3_mAd043_2 CB@3_mAd044_1 CB@3_mAd044_2 CB@3_mAd045_1 CB@3_mAd045_2 CB@3_mAd046_1 CB@3_mAd046_2 CB@3_mAd047_1 CB@3_mAd047_2 CB@3_mAd050_1 CB@3_mAd050_2 CB@3_mAd051_1 CB@3_mAd051_2 CB@3_mAd052_1 CB@3_mAd052_2 CB@3_mAd053_1 CB@3_mAd053_2 CB@3_mAd054_1 CB@3_mAd054_2 CB@3_mAd055_1 CB@3_mAd055_2 CB@3_mAd056_1 CB@3_mAd056_2 CB@3_mAd057_1 CB@3_mAd057_2 CB@3_mAd060_1 CB@3_mAd060_2 CB@3_mAd066_1 
+CB@3_mAd066_2 CB@3_mAd067_1 CB@3_mAd067_2 CB@3_mAd100_1 CB@3_mAd100_2 CB@3_mAd101_1 CB@3_mAd101_2 CB@3_mAd102_1 CB@3_mAd102_2 CB@3_mAd110_1 CB@3_mAd110_2 CB@3_mAd111_1 CB@3_mAd111_2 CB@3_mAd112_1 CB@3_mAd112_2 CB@3_mAd113_1 CB@3_mAd113_2 CB@3_mAd114_1 CB@3_mAd114_2 CB@3_mAd115_1 CB@3_mAd115_2 CB@3_mAd116_1 CB@3_mAd116_2 CB@3_mAd117_1 CB@3_mAd117_2 CB@3_mAd120_1 CB@3_mAd120_2 CB@3_mAd121_1 CB@3_mAd121_2 CB@3_mAd122_1 CB@3_mAd122_2 CB@3_mAd123_1 CB@3_mAd123_2 CB@3_mAd124_1 CB@3_mAd124_2 CB@3_mAd125_1 
+CB@3_mAd125_2 CB@3_mAd126_1 CB@3_mAd126_2 CB@3_mAd127_1 CB@3_mAd127_2 CB@3_mAd130_1 CB@3_mAd130_2 CB@3_mAd131_1 CB@3_mAd131_2 CB@3_mAd132_1 CB@3_mAd132_2 CB@3_mAd133_1 CB@3_mAd133_2 CB@3_mAd134_1 CB@3_mAd134_2 CB@3_mAd135_1 CB@3_mAd135_2 CB@3_mAd136_1 CB@3_mAd136_2 CB@3_mAd137_1 CB@3_mAd137_2 CB@3_mAd140_1 CB@3_mAd140_2 CB@3_mAd141_1 CB@3_mAd141_2 CB@3_mAd142_1 CB@3_mAd142_2 CB@3_mAd143_1 CB@3_mAd143_2 CB@3_mAd144_1 CB@3_mAd144_2 CB@3_mAd145_1 CB@3_mAd145_2 CB@3_mAd146_1 CB@3_mAd146_2 CB@3_mAd147_1 
+CB@3_mAd147_2 CB@3_mAd150_1 CB@3_mAd150_2 CB@3_mAd151_1 CB@3_mAd151_2 CB@3_mAd152_1 CB@3_mAd152_2 CB@3_mAd153_1 CB@3_mAd153_2 CB@3_mAd154_1 CB@3_mAd154_2 CB@3_mAd155_1 CB@3_mAd155_2 CB@3_mAd156_1 CB@3_mAd156_2 CB@3_mAd157_1 CB@3_mAd157_2 CB@3_mAd160_1 CB@3_mAd160_2 CB@3_mAd161_1 CB@3_mAd161_2 CB@3_mAd162_1 CB@3_mAd162_2 CB@3_mAd163_1 CB@3_mAd163_2 CB@3_mAd164_1 CB@3_mAd164_2 CB@3_mAd165_1 CB@3_mAd165_2 CB@3_mAd166_1 CB@3_mAd166_2 CB@3_mAd167_1 CB@3_mAd167_2 CB@3_mAd170_1 CB@3_mAd170_2 CB@3_mAd171_1 
+CB@3_mAd171_2 CB@3_mAd172_1 CB@3_mAd172_2 CB@3_mAd173_1 CB@3_mAd173_2 CB@3_mAd175_1 CB@3_mAd175_2 CB@3_mAd176_1 CB@3_mAd176_2 CB@3_mAd177_1 CB@3_mAd177_2 CB@3_mAd200_1 CB@3_mAd200_2 CB@3_mAd201_1 CB@3_mAd201_2 CB@3_mAd202_1 CB@3_mAd202_2 CB@3_mAd204_1 CB@3_mAd204_2 CB@3_mAd205_1 CB@3_mAd205_2 CB@3_mAd206_1 CB@3_mAd206_2 CB@3_mAd207_1 CB@3_mAd207_2 CB@3_mAd210_1 CB@3_mAd210_2 CB@3_mAd211_1 CB@3_mAd211_2 CB@3_mAd212_1 CB@3_mAd212_2 CB@3_mAd213_1 CB@3_mAd213_2 CB@3_mAd214_1 CB@3_mAd214_2 CB@3_mAd215_1 
+CB@3_mAd215_2 CB@3_mAd216_1 CB@3_mAd216_2 CB@3_mAd217_1 CB@3_mAd217_2 CB@3_mAd220_1 CB@3_mAd220_2 CB@3_mAd221_1 CB@3_mAd221_2 CB@3_mAd222_1 CB@3_mAd222_2 CB@3_mAd223_1 CB@3_mAd223_2 CB@3_mAd224_1 CB@3_mAd224_2 CB@3_mAd225_1 CB@3_mAd225_2 CB@3_mAd226_1 CB@3_mAd226_2 CB@3_mAd227_1 CB@3_mAd227_2 CB@3_mAd230_1 CB@3_mAd230_2 CB@3_mAd231_1 CB@3_mAd231_2 CB@3_mAd232_1 CB@3_mAd232_2 CB@3_mAd233_1 CB@3_mAd233_2 CB@3_mAd234_1 CB@3_mAd234_2 CB@3_mAd235_1 CB@3_mAd235_2 CB@3_mAd236_1 CB@3_mAd236_2 CB@3_mAd237_1 
+CB@3_mAd237_2 CB@3_mAd240_1 CB@3_mAd240_2 CB@3_mAd241_1 CB@3_mAd241_2 CB@3_mAd242_1 CB@3_mAd242_2 CB@3_mAd243_1 CB@3_mAd243_2 CB@3_mAd244_1 CB@3_mAd244_2 CB@3_mAd245_1 CB@3_mAd245_2 CB@3_mAd246_1 CB@3_mAd246_2 CB@3_mAd247_1 CB@3_mAd247_2 CB@3_mAd250_1 CB@3_mAd250_2 CB@3_mAd251_1 CB@3_mAd251_2 CB@3_mAd252_1 CB@3_mAd252_2 CB@3_mAd253_1 CB@3_mAd253_2 CB@3_mAd254_1 CB@3_mAd254_2 CB@3_mAd255_1 CB@3_mAd255_2 CB@3_mAd256_1 CB@3_mAd256_2 CB@3_mAd257_1 CB@3_mAd257_2 CB@3_mAd260_1 CB@3_mAd260_2 CB@3_mAd261_1 
+CB@3_mAd261_2 CB@3_mAd262_1 CB@3_mAd262_2 CB@3_mAd263_1 CB@3_mAd263_2 CB@3_mAd264_1 CB@3_mAd264_2 CB@3_mAd265_1 CB@3_mAd265_2 CB@3_mAd266_1 CB@3_mAd266_2 CB@3_mAd267_1 CB@3_mAd267_2 CB@3_mAd275_1 CB@3_mAd275_2 CB@3_mAd276_1 CB@3_mAd276_2 CB@3_mAd277_1 CB@3_mAd277_2 CB@3_mAd300_1 CB@3_mAd300_2 CB@3_mAd310_1 CB@3_mAd310_2 CB@3_mAd311_1 CB@3_mAd311_2 CB@3_mAd317_1 CB@3_mAd317_2 CB@3_mAd320_1 CB@3_mAd320_2 CB@3_mAd321_1 CB@3_mAd321_2 CB@3_mAd322_1 CB@3_mAd322_2 CB@3_mAd323_1 CB@3_mAd323_2 CB@3_mAd324_1 
+CB@3_mAd324_2 CB@3_mAd325_1 CB@3_mAd325_2 CB@3_mAd326_1 CB@3_mAd326_2 CB@3_mAd327_1 CB@3_mAd327_2 CB@3_mAd330_1 CB@3_mAd330_2 CB@3_mAd331_1 CB@3_mAd331_2 CB@3_mAd332_1 CB@3_mAd332_2 CB@3_mAd333_1 CB@3_mAd333_2 CB@3_mAd334_1 CB@3_mAd334_2 CB@3_mAd335_1 CB@3_mAd335_2 CB@3_mAd336_1 CB@3_mAd336_2 CB@3_mAd337_1 CB@3_mAd337_2 CB@3_mAd340_1 CB@3_mAd340_2 CB@3_mAd341_1 CB@3_mAd341_2 CB@3_mAd342_1 CB@3_mAd342_2 CB@3_mAd343_1 CB@3_mAd343_2 CB@3_mAd344_1 CB@3_mAd344_2 CB@3_mAd345_1 CB@3_mAd345_2 CB@3_mAd346_1 
+CB@3_mAd346_2 CB@3_mAd347_1 CB@3_mAd347_2 CB@3_mAd350_1 CB@3_mAd350_2 CB@3_mAd351_1 CB@3_mAd351_2 CB@3_mAd352_1 CB@3_mAd352_2 CB@3_mAd353_1 CB@3_mAd353_2 CB@3_mAd354_1 CB@3_mAd354_2 CB@3_mAd355_1 CB@3_mAd355_2 CB@3_mAd356_1 CB@3_mAd356_2 CB@3_mAd357_1 CB@3_mAd357_2 CB@3_mAd360_1 CB@3_mAd360_2 CB@3_mAd361_1 CB@3_mAd361_2 CB@3_mAd362_1 CB@3_mAd362_2 CB@3_mAd363_1 CB@3_mAd363_2 CB@3_mAd364_1 CB@3_mAd364_2 CB@3_mAd365_1 CB@3_mAd365_2 CB@3_mAd366_1 CB@3_mAd366_2 CB@3_mAd367_1 CB@3_mAd367_2 CB@3_mAd371_1 
+CB@3_mAd371_2 CB@3_mAd372_1 CB@3_mAd372_2 CB@3_mAd373_1 CB@3_mAd373_2 CB@3_mAd374_1 CB@3_mAd374_2 CB@3_mAd375_1 CB@3_mAd375_2 CB@3_mAd376_1 CB@3_mAd376_2 CB@3_mAd377_1 CB@3_mAd377_2 CB@3_mAd400_1 CB@3_mAd400_2 CB@3_mAd401_1 CB@3_mAd401_2 CB@3_mAd402_1 CB@3_mAd402_2 CB@3_mAd403_1 CB@3_mAd403_2 CB@3_mAd404_1 CB@3_mAd404_2 CB@3_mAd405_1 CB@3_mAd405_2 CB@3_mAd406_1 CB@3_mAd406_2 CB@3_mAd407_1 CB@3_mAd407_2 CB@3_mAd410_1 CB@3_mAd410_2 CB@3_mAd411_1 CB@3_mAd411_2 CB@3_mAd412_1 CB@3_mAd412_2 CB@3_mAd413_1 
+CB@3_mAd413_2 CB@3_mAd414_1 CB@3_mAd414_2 CB@3_mAd415_1 CB@3_mAd415_2 CB@3_mAd416_1 CB@3_mAd416_2 CB@3_mAd417_1 CB@3_mAd417_2 CB@3_mAd420_1 CB@3_mAd420_2 CB@3_mAd421_1 CB@3_mAd421_2 CB@3_mAd422_1 CB@3_mAd422_2 CB@3_mAd423_1 CB@3_mAd423_2 CB@3_mAd424_1 CB@3_mAd424_2 CB@3_mAd425_1 CB@3_mAd425_2 CB@3_mAd426_1 CB@3_mAd426_2 CB@3_mAd427_1 CB@3_mAd427_2 CB@3_mAd430_1 CB@3_mAd430_2 CB@3_mAd431_1 CB@3_mAd431_2 CB@3_mAd432_1 CB@3_mAd432_2 CB@3_mAd433_1 CB@3_mAd433_2 CB@3_mAd434_1 CB@3_mAd434_2 CB@3_mAd435_1 
+CB@3_mAd435_2 CB@3_mAd436_1 CB@3_mAd436_2 CB@3_mAd437_1 CB@3_mAd437_2 CB@3_mAd440_1 CB@3_mAd440_2 CB@3_mAd441_1 CB@3_mAd441_2 CB@3_mAd442_1 CB@3_mAd442_2 CB@3_mAd443_1 CB@3_mAd443_2 CB@3_mAd444_1 CB@3_mAd444_2 CB@3_mAd445_1 CB@3_mAd445_2 CB@3_mAd446_1 CB@3_mAd446_2 CB@3_mAd447_1 CB@3_mAd447_2 CB@3_mAd450_1 CB@3_mAd450_2 CB@3_mAd451_1 CB@3_mAd451_2 CB@3_mAd452_1 CB@3_mAd452_2 CB@3_mAd453_1 CB@3_mAd453_2 CB@3_mAd454_1 CB@3_mAd454_2 CB@3_mAd455_1 CB@3_mAd455_2 CB@3_mAd456_1 CB@3_mAd456_2 CB@3_mAd457_1 
+CB@3_mAd457_2 CB@3_mAd460_1 CB@3_mAd460_2 CB@3_mAd466_1 CB@3_mAd466_2 CB@3_mAd467_1 CB@3_mAd467_2 CB@3_mAd500_1 CB@3_mAd500_2 CB@3_mAd501_1 CB@3_mAd501_2 CB@3_mAd502_1 CB@3_mAd502_2 CB@3_mAd508_1 CB@3_mAd508_2 CB@3_mAd509_1 CB@3_mAd509_2 CB@3_mAd512_1 CB@3_mAd512_2 CB@3_mAd513_1 CB@3_mAd513_2 CB@3_mAd514_1 CB@3_mAd514_2 CB@3_mAd515_1 CB@3_mAd515_2 CB@3_mAd516_1 CB@3_mAd516_2 CB@3_mAd517_1 CB@3_mAd517_2 CB@3_mAd520_1 CB@3_mAd520_2 CB@3_mAd521_1 CB@3_mAd521_2 CB@3_mAd522_1 CB@3_mAd522_2 CB@3_mAd523_1 
+CB@3_mAd523_2 CB@3_mAd524_1 CB@3_mAd524_2 CB@3_mAd525_1 CB@3_mAd525_2 CB@3_mAd526_1 CB@3_mAd526_2 CB@3_mAd527_1 CB@3_mAd527_2 CB@3_mAd530_1 CB@3_mAd530_2 CB@3_mAd531_1 CB@3_mAd531_2 CB@3_mAd532_1 CB@3_mAd532_2 CB@3_mAd533_1 CB@3_mAd533_2 CB@3_mAd534_1 CB@3_mAd534_2 CB@3_mAd535_1 CB@3_mAd535_2 CB@3_mAd536_1 CB@3_mAd536_2 CB@3_mAd537_1 CB@3_mAd537_2 CB@3_mAd540_1 CB@3_mAd540_2 CB@3_mAd541_1 CB@3_mAd541_2 CB@3_mAd542_1 CB@3_mAd542_2 CB@3_mAd543_1 CB@3_mAd543_2 CB@3_mAd544_1 CB@3_mAd544_2 CB@3_mAd545_1 
+CB@3_mAd545_2 CB@3_mAd546_1 CB@3_mAd546_2 CB@3_mAd547_1 CB@3_mAd547_2 CB@3_mAd550_1 CB@3_mAd550_2 CB@3_mAd551_1 CB@3_mAd551_2 CB@3_mAd552_1 CB@3_mAd552_2 CB@3_mAd553_1 CB@3_mAd553_2 CB@3_mAd554_1 CB@3_mAd554_2 CB@3_mAd555_1 CB@3_mAd555_2 CB@3_mAd556_1 CB@3_mAd556_2 CB@3_mAd557_1 CB@3_mAd557_2 CB@3_mAd560_1 CB@3_mAd560_2 CB@3_mAd561_1 CB@3_mAd561_2 CB@3_mAd562_1 CB@3_mAd562_2 CB@3_mAd563_1 CB@3_mAd563_2 CB@3_mAd564_1 CB@3_mAd564_2 CB@3_mAd565_1 CB@3_mAd565_2 CB@3_mAd566_1 CB@3_mAd566_2 CB@3_mAd567_1 
+CB@3_mAd567_2 CB@3_mAd570_1 CB@3_mAd570_2 CB@3_mAd571_1 CB@3_mAd571_2 CB@3_mAd572_1 CB@3_mAd572_2 CB@3_mAd573_1 CB@3_mAd573_2 CB@3_mAd575_1 CB@3_mAd575_2 CB@3_mAd576_1 CB@3_mAd576_2 CB@3_mAd577_1 CB@3_mAd577_2 CB@3_mAd600_1 CB@3_mAd600_2 CB@3_mAd601_1 CB@3_mAd601_2 CB@3_mAd602_1 CB@3_mAd602_2 CB@3_mAd604_1 CB@3_mAd604_2 CB@3_mAd605_1 CB@3_mAd605_2 CB@3_mAd606_1 CB@3_mAd606_2 CB@3_mAd607_1 CB@3_mAd607_2 CB@3_mAd610_1 CB@3_mAd610_2 CB@3_mAd611_1 CB@3_mAd611_2 CB@3_mAd612_1 CB@3_mAd612_2 CB@3_mAd613_1 
+CB@3_mAd613_2 CB@3_mAd614_1 CB@3_mAd614_2 CB@3_mAd615_1 CB@3_mAd615_2 CB@3_mAd616_1 CB@3_mAd616_2 CB@3_mAd617_1 CB@3_mAd617_2 CB@3_mAd620_1 CB@3_mAd620_2 CB@3_mAd621_1 CB@3_mAd621_2 CB@3_mAd622_1 CB@3_mAd622_2 CB@3_mAd623_1 CB@3_mAd623_2 CB@3_mAd624_1 CB@3_mAd624_2 CB@3_mAd625_1 CB@3_mAd625_2 CB@3_mAd626_1 CB@3_mAd626_2 CB@3_mAd627_1 CB@3_mAd627_2 CB@3_mAd630_1 CB@3_mAd630_2 CB@3_mAd631_1 CB@3_mAd631_2 CB@3_mAd632_1 CB@3_mAd632_2 CB@3_mAd633_1 CB@3_mAd633_2 CB@3_mAd634_1 CB@3_mAd634_2 CB@3_mAd635_1 
+CB@3_mAd635_2 CB@3_mAd636_1 CB@3_mAd636_2 CB@3_mAd637_1 CB@3_mAd637_2 CB@3_mAd640_1 CB@3_mAd640_2 CB@3_mAd641_1 CB@3_mAd641_2 CB@3_mAd642_1 CB@3_mAd642_2 CB@3_mAd643_1 CB@3_mAd643_2 CB@3_mAd644_1 CB@3_mAd644_2 CB@3_mAd645_1 CB@3_mAd645_2 CB@3_mAd646_1 CB@3_mAd646_2 CB@3_mAd647_1 CB@3_mAd647_2 CB@3_mAd650_1 CB@3_mAd650_2 CB@3_mAd651_1 CB@3_mAd651_2 CB@3_mAd652_1 CB@3_mAd652_2 CB@3_mAd653_1 CB@3_mAd653_2 CB@3_mAd654_1 CB@3_mAd654_2 CB@3_mAd655_1 CB@3_mAd655_2 CB@3_mAd656_1 CB@3_mAd656_2 CB@3_mAd657_1 
+CB@3_mAd657_2 CB@3_mAd660_1 CB@3_mAd660_2 CB@3_mAd661_1 CB@3_mAd661_2 CB@3_mAd662_1 CB@3_mAd662_2 CB@3_mAd663_1 CB@3_mAd663_2 CB@3_mAd664_1 CB@3_mAd664_2 CB@3_mAd665_1 CB@3_mAd665_2 CB@3_mAd666_1 CB@3_mAd666_2 CB@3_mAd667_1 CB@3_mAd667_2 CB@3_mAd675_1 CB@3_mAd675_2 CB@3_mAd676_1 CB@3_mAd676_2 CB@3_mAd677_1 CB@3_mAd677_2 CB@3_mAd700_1 CB@3_mAd700_2 CB@3_mAd710_1 CB@3_mAd710_2 CB@3_mAd711_1 CB@3_mAd711_2 CB@3_mAd717_1 CB@3_mAd717_2 CB@3_mAd720_1 CB@3_mAd720_2 CB@3_mAd721_1 CB@3_mAd721_2 CB@3_mAd722_1 
+CB@3_mAd722_2 CB@3_mAd723_1 CB@3_mAd723_2 CB@3_mAd724_1 CB@3_mAd724_2 CB@3_mAd725_1 CB@3_mAd725_2 CB@3_mAd726_1 CB@3_mAd726_2 CB@3_mAd727_1 CB@3_mAd727_2 CB@3_mAd730_1 CB@3_mAd730_2 CB@3_mAd731_1 CB@3_mAd731_2 CB@3_mAd732_1 CB@3_mAd732_2 CB@3_mAd733_1 CB@3_mAd733_2 CB@3_mAd734_1 CB@3_mAd734_2 CB@3_mAd735_1 CB@3_mAd735_2 CB@3_mAd736_1 CB@3_mAd736_2 CB@3_mAd737_1 CB@3_mAd737_2 CB@3_mAd740_1 CB@3_mAd740_2 CB@3_mAd741_1 CB@3_mAd741_2 CB@3_mAd742_1 CB@3_mAd742_2 CB@3_mAd743_1 CB@3_mAd743_2 CB@3_mAd744_1 
+CB@3_mAd744_2 CB@3_mAd745_1 CB@3_mAd745_2 CB@3_mAd746_1 CB@3_mAd746_2 CB@3_mAd747_1 CB@3_mAd747_2 CB@3_mAd750_1 CB@3_mAd750_2 CB@3_mAd751_1 CB@3_mAd751_2 CB@3_mAd752_1 CB@3_mAd752_2 CB@3_mAd753_1 CB@3_mAd753_2 CB@3_mAd754_1 CB@3_mAd754_2 CB@3_mAd755_1 CB@3_mAd755_2 CB@3_mAd756_1 CB@3_mAd756_2 CB@3_mAd757_1 CB@3_mAd757_2 CB@3_mAd760_1 CB@3_mAd760_2 CB@3_mAd761_1 CB@3_mAd761_2 CB@3_mAd762_1 CB@3_mAd762_2 CB@3_mAd763_1 CB@3_mAd763_2 CB@3_mAd764_1 CB@3_mAd764_2 CB@3_mAd765_1 CB@3_mAd765_2 CB@3_mAd766_1 
+CB@3_mAd766_2 CB@3_mAd767_1 CB@3_mAd767_2 CB@3_mAd771_1 CB@3_mAd771_2 CB@3_mAd772_1 CB@3_mAd772_2 CB@3_mAd773_1 CB@3_mAd773_2 CB@3_mAd774_1 CB@3_mAd774_2 CB@3_mAd775_1 CB@3_mAd775_2 CB@3_mAd776_1 CB@3_mAd776_2 CB@3_mAd777_1 CB@3_mAd777_2 CB@3_X0 CB@3_X1 CB@3_X10 CB@3_X11 CB@3_X12 CB@3_X13 CB@3_X2 CB@3_X3 CB@3_X4 CB@3_X5 CB@3_X6 CB@3_X7 CB@3_X8 CB@3_X9 CB@3_Y1 CB@3_Y10 CB@3_Y11 CB@3_Y12 CB@3_Y2 CB@3_Y3 CB@3_Y4 CB@3_Y5 CB@3_Y6 CB@3_Y7 CB@3_Y8 CB@3_Y9 CB@3_Z1 CB@3_Z10 CB@3_Z11 CB@3_Z12 CB@3_Z2 CB@3_Z3 CB@3_Z4 
+CB@3_Z5 CB@3_Z6 CB@3_Z7 CB@3_Z8 CB@3_Z9 _5400TP094__CB
XCB@4 CB@4_K0 CB@4_K1 CB@4_K10 CB@4_K11 CB@4_K12 CB@4_K13 CB@4_K2 CB@4_K3 CB@4_K4 CB@4_K5 CB@4_K6 CB@4_K7 CB@4_K8 CB@4_K9 CB@4_mAd000_1 CB@4_mAd000_2 CB@4_mAd001_1 CB@4_mAd001_2 CB@4_mAd002_1 CB@4_mAd002_2 CB@4_mAd003_1 CB@4_mAd003_2 CB@4_mAd004_1 CB@4_mAd004_2 CB@4_mAd005_1 CB@4_mAd005_2 CB@4_mAd006_1 CB@4_mAd006_2 CB@4_mAd007_1 CB@4_mAd007_2 CB@4_mAd010_1 CB@4_mAd010_2 CB@4_mAd011_1 CB@4_mAd011_2 CB@4_mAd012_1 CB@4_mAd012_2 CB@4_mAd013_1 CB@4_mAd013_2 CB@4_mAd014_1 CB@4_mAd014_2 CB@4_mAd015_1 
+CB@4_mAd015_2 CB@4_mAd016_1 CB@4_mAd016_2 CB@4_mAd017_1 CB@4_mAd017_2 CB@4_mAd020_1 CB@4_mAd020_2 CB@4_mAd021_1 CB@4_mAd021_2 CB@4_mAd022_1 CB@4_mAd022_2 CB@4_mAd023_1 CB@4_mAd023_2 CB@4_mAd024_1 CB@4_mAd024_2 CB@4_mAd025_1 CB@4_mAd025_2 CB@4_mAd026_1 CB@4_mAd026_2 CB@4_mAd027_1 CB@4_mAd027_2 CB@4_mAd030_1 CB@4_mAd030_2 CB@4_mAd031_1 CB@4_mAd031_2 CB@4_mAd032_1 CB@4_mAd032_2 CB@4_mAd033_1 CB@4_mAd033_2 CB@4_mAd034_1 CB@4_mAd034_2 CB@4_mAd035_1 CB@4_mAd035_2 CB@4_mAd036_1 CB@4_mAd036_2 CB@4_mAd037_1 
+CB@4_mAd037_2 CB@4_mAd040_1 CB@4_mAd040_2 CB@4_mAd041_1 CB@4_mAd041_2 CB@4_mAd042_1 CB@4_mAd042_2 CB@4_mAd043_1 CB@4_mAd043_2 CB@4_mAd044_1 CB@4_mAd044_2 CB@4_mAd045_1 CB@4_mAd045_2 CB@4_mAd046_1 CB@4_mAd046_2 CB@4_mAd047_1 CB@4_mAd047_2 CB@4_mAd050_1 CB@4_mAd050_2 CB@4_mAd051_1 CB@4_mAd051_2 CB@4_mAd052_1 CB@4_mAd052_2 CB@4_mAd053_1 CB@4_mAd053_2 CB@4_mAd054_1 CB@4_mAd054_2 CB@4_mAd055_1 CB@4_mAd055_2 CB@4_mAd056_1 CB@4_mAd056_2 CB@4_mAd057_1 CB@4_mAd057_2 CB@4_mAd060_1 CB@4_mAd060_2 CB@4_mAd066_1 
+CB@4_mAd066_2 CB@4_mAd067_1 CB@4_mAd067_2 CB@4_mAd100_1 CB@4_mAd100_2 CB@4_mAd101_1 CB@4_mAd101_2 CB@4_mAd102_1 CB@4_mAd102_2 CB@4_mAd110_1 CB@4_mAd110_2 CB@4_mAd111_1 CB@4_mAd111_2 CB@4_mAd112_1 CB@4_mAd112_2 CB@4_mAd113_1 CB@4_mAd113_2 CB@4_mAd114_1 CB@4_mAd114_2 CB@4_mAd115_1 CB@4_mAd115_2 CB@4_mAd116_1 CB@4_mAd116_2 CB@4_mAd117_1 CB@4_mAd117_2 CB@4_mAd120_1 CB@4_mAd120_2 CB@4_mAd121_1 CB@4_mAd121_2 CB@4_mAd122_1 CB@4_mAd122_2 CB@4_mAd123_1 CB@4_mAd123_2 CB@4_mAd124_1 CB@4_mAd124_2 CB@4_mAd125_1 
+CB@4_mAd125_2 CB@4_mAd126_1 CB@4_mAd126_2 CB@4_mAd127_1 CB@4_mAd127_2 CB@4_mAd130_1 CB@4_mAd130_2 CB@4_mAd131_1 CB@4_mAd131_2 CB@4_mAd132_1 CB@4_mAd132_2 CB@4_mAd133_1 CB@4_mAd133_2 CB@4_mAd134_1 CB@4_mAd134_2 CB@4_mAd135_1 CB@4_mAd135_2 CB@4_mAd136_1 CB@4_mAd136_2 CB@4_mAd137_1 CB@4_mAd137_2 CB@4_mAd140_1 CB@4_mAd140_2 CB@4_mAd141_1 CB@4_mAd141_2 CB@4_mAd142_1 CB@4_mAd142_2 CB@4_mAd143_1 CB@4_mAd143_2 CB@4_mAd144_1 CB@4_mAd144_2 CB@4_mAd145_1 CB@4_mAd145_2 CB@4_mAd146_1 CB@4_mAd146_2 CB@4_mAd147_1 
+CB@4_mAd147_2 CB@4_mAd150_1 CB@4_mAd150_2 CB@4_mAd151_1 CB@4_mAd151_2 CB@4_mAd152_1 CB@4_mAd152_2 CB@4_mAd153_1 CB@4_mAd153_2 CB@4_mAd154_1 CB@4_mAd154_2 CB@4_mAd155_1 CB@4_mAd155_2 CB@4_mAd156_1 CB@4_mAd156_2 CB@4_mAd157_1 CB@4_mAd157_2 CB@4_mAd160_1 CB@4_mAd160_2 CB@4_mAd161_1 CB@4_mAd161_2 CB@4_mAd162_1 CB@4_mAd162_2 CB@4_mAd163_1 CB@4_mAd163_2 CB@4_mAd164_1 CB@4_mAd164_2 CB@4_mAd165_1 CB@4_mAd165_2 CB@4_mAd166_1 CB@4_mAd166_2 CB@4_mAd167_1 CB@4_mAd167_2 CB@4_mAd170_1 CB@4_mAd170_2 CB@4_mAd171_1 
+CB@4_mAd171_2 CB@4_mAd172_1 CB@4_mAd172_2 CB@4_mAd173_1 CB@4_mAd173_2 CB@4_mAd175_1 CB@4_mAd175_2 CB@4_mAd176_1 CB@4_mAd176_2 CB@4_mAd177_1 CB@4_mAd177_2 CB@4_mAd200_1 CB@4_mAd200_2 CB@4_mAd201_1 CB@4_mAd201_2 CB@4_mAd202_1 CB@4_mAd202_2 CB@4_mAd204_1 CB@4_mAd204_2 CB@4_mAd205_1 CB@4_mAd205_2 CB@4_mAd206_1 CB@4_mAd206_2 CB@4_mAd207_1 CB@4_mAd207_2 CB@4_mAd210_1 CB@4_mAd210_2 CB@4_mAd211_1 CB@4_mAd211_2 CB@4_mAd212_1 CB@4_mAd212_2 CB@4_mAd213_1 CB@4_mAd213_2 CB@4_mAd214_1 CB@4_mAd214_2 CB@4_mAd215_1 
+CB@4_mAd215_2 CB@4_mAd216_1 CB@4_mAd216_2 CB@4_mAd217_1 CB@4_mAd217_2 CB@4_mAd220_1 CB@4_mAd220_2 CB@4_mAd221_1 CB@4_mAd221_2 CB@4_mAd222_1 CB@4_mAd222_2 CB@4_mAd223_1 CB@4_mAd223_2 CB@4_mAd224_1 CB@4_mAd224_2 CB@4_mAd225_1 CB@4_mAd225_2 CB@4_mAd226_1 CB@4_mAd226_2 CB@4_mAd227_1 CB@4_mAd227_2 CB@4_mAd230_1 CB@4_mAd230_2 CB@4_mAd231_1 CB@4_mAd231_2 CB@4_mAd232_1 CB@4_mAd232_2 CB@4_mAd233_1 CB@4_mAd233_2 CB@4_mAd234_1 CB@4_mAd234_2 CB@4_mAd235_1 CB@4_mAd235_2 CB@4_mAd236_1 CB@4_mAd236_2 CB@4_mAd237_1 
+CB@4_mAd237_2 CB@4_mAd240_1 CB@4_mAd240_2 CB@4_mAd241_1 CB@4_mAd241_2 CB@4_mAd242_1 CB@4_mAd242_2 CB@4_mAd243_1 CB@4_mAd243_2 CB@4_mAd244_1 CB@4_mAd244_2 CB@4_mAd245_1 CB@4_mAd245_2 CB@4_mAd246_1 CB@4_mAd246_2 CB@4_mAd247_1 CB@4_mAd247_2 CB@4_mAd250_1 CB@4_mAd250_2 CB@4_mAd251_1 CB@4_mAd251_2 CB@4_mAd252_1 CB@4_mAd252_2 CB@4_mAd253_1 CB@4_mAd253_2 CB@4_mAd254_1 CB@4_mAd254_2 CB@4_mAd255_1 CB@4_mAd255_2 CB@4_mAd256_1 CB@4_mAd256_2 CB@4_mAd257_1 CB@4_mAd257_2 CB@4_mAd260_1 CB@4_mAd260_2 CB@4_mAd261_1 
+CB@4_mAd261_2 CB@4_mAd262_1 CB@4_mAd262_2 CB@4_mAd263_1 CB@4_mAd263_2 CB@4_mAd264_1 CB@4_mAd264_2 CB@4_mAd265_1 CB@4_mAd265_2 CB@4_mAd266_1 CB@4_mAd266_2 CB@4_mAd267_1 CB@4_mAd267_2 CB@4_mAd275_1 CB@4_mAd275_2 CB@4_mAd276_1 CB@4_mAd276_2 CB@4_mAd277_1 CB@4_mAd277_2 CB@4_mAd300_1 CB@4_mAd300_2 CB@4_mAd310_1 CB@4_mAd310_2 CB@4_mAd311_1 CB@4_mAd311_2 CB@4_mAd317_1 CB@4_mAd317_2 CB@4_mAd320_1 CB@4_mAd320_2 CB@4_mAd321_1 CB@4_mAd321_2 CB@4_mAd322_1 CB@4_mAd322_2 CB@4_mAd323_1 CB@4_mAd323_2 CB@4_mAd324_1 
+CB@4_mAd324_2 CB@4_mAd325_1 CB@4_mAd325_2 CB@4_mAd326_1 CB@4_mAd326_2 CB@4_mAd327_1 CB@4_mAd327_2 CB@4_mAd330_1 CB@4_mAd330_2 CB@4_mAd331_1 CB@4_mAd331_2 CB@4_mAd332_1 CB@4_mAd332_2 CB@4_mAd333_1 CB@4_mAd333_2 CB@4_mAd334_1 CB@4_mAd334_2 CB@4_mAd335_1 CB@4_mAd335_2 CB@4_mAd336_1 CB@4_mAd336_2 CB@4_mAd337_1 CB@4_mAd337_2 CB@4_mAd340_1 CB@4_mAd340_2 CB@4_mAd341_1 CB@4_mAd341_2 CB@4_mAd342_1 CB@4_mAd342_2 CB@4_mAd343_1 CB@4_mAd343_2 CB@4_mAd344_1 CB@4_mAd344_2 CB@4_mAd345_1 CB@4_mAd345_2 CB@4_mAd346_1 
+CB@4_mAd346_2 CB@4_mAd347_1 CB@4_mAd347_2 CB@4_mAd350_1 CB@4_mAd350_2 CB@4_mAd351_1 CB@4_mAd351_2 CB@4_mAd352_1 CB@4_mAd352_2 CB@4_mAd353_1 CB@4_mAd353_2 CB@4_mAd354_1 CB@4_mAd354_2 CB@4_mAd355_1 CB@4_mAd355_2 CB@4_mAd356_1 CB@4_mAd356_2 CB@4_mAd357_1 CB@4_mAd357_2 CB@4_mAd360_1 CB@4_mAd360_2 CB@4_mAd361_1 CB@4_mAd361_2 CB@4_mAd362_1 CB@4_mAd362_2 CB@4_mAd363_1 CB@4_mAd363_2 CB@4_mAd364_1 CB@4_mAd364_2 CB@4_mAd365_1 CB@4_mAd365_2 CB@4_mAd366_1 CB@4_mAd366_2 CB@4_mAd367_1 CB@4_mAd367_2 CB@4_mAd371_1 
+CB@4_mAd371_2 CB@4_mAd372_1 CB@4_mAd372_2 CB@4_mAd373_1 CB@4_mAd373_2 CB@4_mAd374_1 CB@4_mAd374_2 CB@4_mAd375_1 CB@4_mAd375_2 CB@4_mAd376_1 CB@4_mAd376_2 CB@4_mAd377_1 CB@4_mAd377_2 CB@4_mAd400_1 CB@4_mAd400_2 CB@4_mAd401_1 CB@4_mAd401_2 CB@4_mAd402_1 CB@4_mAd402_2 CB@4_mAd403_1 CB@4_mAd403_2 CB@4_mAd404_1 CB@4_mAd404_2 CB@4_mAd405_1 CB@4_mAd405_2 CB@4_mAd406_1 CB@4_mAd406_2 CB@4_mAd407_1 CB@4_mAd407_2 CB@4_mAd410_1 CB@4_mAd410_2 CB@4_mAd411_1 CB@4_mAd411_2 CB@4_mAd412_1 CB@4_mAd412_2 CB@4_mAd413_1 
+CB@4_mAd413_2 CB@4_mAd414_1 CB@4_mAd414_2 CB@4_mAd415_1 CB@4_mAd415_2 CB@4_mAd416_1 CB@4_mAd416_2 CB@4_mAd417_1 CB@4_mAd417_2 CB@4_mAd420_1 CB@4_mAd420_2 CB@4_mAd421_1 CB@4_mAd421_2 CB@4_mAd422_1 CB@4_mAd422_2 CB@4_mAd423_1 CB@4_mAd423_2 CB@4_mAd424_1 CB@4_mAd424_2 CB@4_mAd425_1 CB@4_mAd425_2 CB@4_mAd426_1 CB@4_mAd426_2 CB@4_mAd427_1 CB@4_mAd427_2 CB@4_mAd430_1 CB@4_mAd430_2 CB@4_mAd431_1 CB@4_mAd431_2 CB@4_mAd432_1 CB@4_mAd432_2 CB@4_mAd433_1 CB@4_mAd433_2 CB@4_mAd434_1 CB@4_mAd434_2 CB@4_mAd435_1 
+CB@4_mAd435_2 CB@4_mAd436_1 CB@4_mAd436_2 CB@4_mAd437_1 CB@4_mAd437_2 CB@4_mAd440_1 CB@4_mAd440_2 CB@4_mAd441_1 CB@4_mAd441_2 CB@4_mAd442_1 CB@4_mAd442_2 CB@4_mAd443_1 CB@4_mAd443_2 CB@4_mAd444_1 CB@4_mAd444_2 CB@4_mAd445_1 CB@4_mAd445_2 CB@4_mAd446_1 CB@4_mAd446_2 CB@4_mAd447_1 CB@4_mAd447_2 CB@4_mAd450_1 CB@4_mAd450_2 CB@4_mAd451_1 CB@4_mAd451_2 CB@4_mAd452_1 CB@4_mAd452_2 CB@4_mAd453_1 CB@4_mAd453_2 CB@4_mAd454_1 CB@4_mAd454_2 CB@4_mAd455_1 CB@4_mAd455_2 CB@4_mAd456_1 CB@4_mAd456_2 CB@4_mAd457_1 
+CB@4_mAd457_2 CB@4_mAd460_1 CB@4_mAd460_2 CB@4_mAd466_1 CB@4_mAd466_2 CB@4_mAd467_1 CB@4_mAd467_2 CB@4_mAd500_1 CB@4_mAd500_2 CB@4_mAd501_1 CB@4_mAd501_2 CB@4_mAd502_1 CB@4_mAd502_2 CB@4_mAd508_1 CB@4_mAd508_2 CB@4_mAd509_1 CB@4_mAd509_2 CB@4_mAd512_1 CB@4_mAd512_2 CB@4_mAd513_1 CB@4_mAd513_2 CB@4_mAd514_1 CB@4_mAd514_2 CB@4_mAd515_1 CB@4_mAd515_2 CB@4_mAd516_1 CB@4_mAd516_2 CB@4_mAd517_1 CB@4_mAd517_2 CB@4_mAd520_1 CB@4_mAd520_2 CB@4_mAd521_1 CB@4_mAd521_2 CB@4_mAd522_1 CB@4_mAd522_2 CB@4_mAd523_1 
+CB@4_mAd523_2 CB@4_mAd524_1 CB@4_mAd524_2 CB@4_mAd525_1 CB@4_mAd525_2 CB@4_mAd526_1 CB@4_mAd526_2 CB@4_mAd527_1 CB@4_mAd527_2 CB@4_mAd530_1 CB@4_mAd530_2 CB@4_mAd531_1 CB@4_mAd531_2 CB@4_mAd532_1 CB@4_mAd532_2 CB@4_mAd533_1 CB@4_mAd533_2 CB@4_mAd534_1 CB@4_mAd534_2 CB@4_mAd535_1 CB@4_mAd535_2 CB@4_mAd536_1 CB@4_mAd536_2 CB@4_mAd537_1 CB@4_mAd537_2 CB@4_mAd540_1 CB@4_mAd540_2 CB@4_mAd541_1 CB@4_mAd541_2 CB@4_mAd542_1 CB@4_mAd542_2 CB@4_mAd543_1 CB@4_mAd543_2 CB@4_mAd544_1 CB@4_mAd544_2 CB@4_mAd545_1 
+CB@4_mAd545_2 CB@4_mAd546_1 CB@4_mAd546_2 CB@4_mAd547_1 CB@4_mAd547_2 CB@4_mAd550_1 CB@4_mAd550_2 CB@4_mAd551_1 CB@4_mAd551_2 CB@4_mAd552_1 CB@4_mAd552_2 CB@4_mAd553_1 CB@4_mAd553_2 CB@4_mAd554_1 CB@4_mAd554_2 CB@4_mAd555_1 CB@4_mAd555_2 CB@4_mAd556_1 CB@4_mAd556_2 CB@4_mAd557_1 CB@4_mAd557_2 CB@4_mAd560_1 CB@4_mAd560_2 CB@4_mAd561_1 CB@4_mAd561_2 CB@4_mAd562_1 CB@4_mAd562_2 CB@4_mAd563_1 CB@4_mAd563_2 CB@4_mAd564_1 CB@4_mAd564_2 CB@4_mAd565_1 CB@4_mAd565_2 CB@4_mAd566_1 CB@4_mAd566_2 CB@4_mAd567_1 
+CB@4_mAd567_2 CB@4_mAd570_1 CB@4_mAd570_2 CB@4_mAd571_1 CB@4_mAd571_2 CB@4_mAd572_1 CB@4_mAd572_2 CB@4_mAd573_1 CB@4_mAd573_2 CB@4_mAd575_1 CB@4_mAd575_2 CB@4_mAd576_1 CB@4_mAd576_2 CB@4_mAd577_1 CB@4_mAd577_2 CB@4_mAd600_1 CB@4_mAd600_2 CB@4_mAd601_1 CB@4_mAd601_2 CB@4_mAd602_1 CB@4_mAd602_2 CB@4_mAd604_1 CB@4_mAd604_2 CB@4_mAd605_1 CB@4_mAd605_2 CB@4_mAd606_1 CB@4_mAd606_2 CB@4_mAd607_1 CB@4_mAd607_2 CB@4_mAd610_1 CB@4_mAd610_2 CB@4_mAd611_1 CB@4_mAd611_2 CB@4_mAd612_1 CB@4_mAd612_2 CB@4_mAd613_1 
+CB@4_mAd613_2 CB@4_mAd614_1 CB@4_mAd614_2 CB@4_mAd615_1 CB@4_mAd615_2 CB@4_mAd616_1 CB@4_mAd616_2 CB@4_mAd617_1 CB@4_mAd617_2 CB@4_mAd620_1 CB@4_mAd620_2 CB@4_mAd621_1 CB@4_mAd621_2 CB@4_mAd622_1 CB@4_mAd622_2 CB@4_mAd623_1 CB@4_mAd623_2 CB@4_mAd624_1 CB@4_mAd624_2 CB@4_mAd625_1 CB@4_mAd625_2 CB@4_mAd626_1 CB@4_mAd626_2 CB@4_mAd627_1 CB@4_mAd627_2 CB@4_mAd630_1 CB@4_mAd630_2 CB@4_mAd631_1 CB@4_mAd631_2 CB@4_mAd632_1 CB@4_mAd632_2 CB@4_mAd633_1 CB@4_mAd633_2 CB@4_mAd634_1 CB@4_mAd634_2 CB@4_mAd635_1 
+CB@4_mAd635_2 CB@4_mAd636_1 CB@4_mAd636_2 CB@4_mAd637_1 CB@4_mAd637_2 CB@4_mAd640_1 CB@4_mAd640_2 CB@4_mAd641_1 CB@4_mAd641_2 CB@4_mAd642_1 CB@4_mAd642_2 CB@4_mAd643_1 CB@4_mAd643_2 CB@4_mAd644_1 CB@4_mAd644_2 CB@4_mAd645_1 CB@4_mAd645_2 CB@4_mAd646_1 CB@4_mAd646_2 CB@4_mAd647_1 CB@4_mAd647_2 CB@4_mAd650_1 CB@4_mAd650_2 CB@4_mAd651_1 CB@4_mAd651_2 CB@4_mAd652_1 CB@4_mAd652_2 CB@4_mAd653_1 CB@4_mAd653_2 CB@4_mAd654_1 CB@4_mAd654_2 CB@4_mAd655_1 CB@4_mAd655_2 CB@4_mAd656_1 CB@4_mAd656_2 CB@4_mAd657_1 
+CB@4_mAd657_2 CB@4_mAd660_1 CB@4_mAd660_2 CB@4_mAd661_1 CB@4_mAd661_2 CB@4_mAd662_1 CB@4_mAd662_2 CB@4_mAd663_1 CB@4_mAd663_2 CB@4_mAd664_1 CB@4_mAd664_2 CB@4_mAd665_1 CB@4_mAd665_2 CB@4_mAd666_1 CB@4_mAd666_2 CB@4_mAd667_1 CB@4_mAd667_2 CB@4_mAd675_1 CB@4_mAd675_2 CB@4_mAd676_1 CB@4_mAd676_2 CB@4_mAd677_1 CB@4_mAd677_2 CB@4_mAd700_1 CB@4_mAd700_2 CB@4_mAd710_1 CB@4_mAd710_2 CB@4_mAd711_1 CB@4_mAd711_2 CB@4_mAd717_1 CB@4_mAd717_2 CB@4_mAd720_1 CB@4_mAd720_2 CB@4_mAd721_1 CB@4_mAd721_2 CB@4_mAd722_1 
+CB@4_mAd722_2 CB@4_mAd723_1 CB@4_mAd723_2 CB@4_mAd724_1 CB@4_mAd724_2 CB@4_mAd725_1 CB@4_mAd725_2 CB@4_mAd726_1 CB@4_mAd726_2 CB@4_mAd727_1 CB@4_mAd727_2 CB@4_mAd730_1 CB@4_mAd730_2 CB@4_mAd731_1 CB@4_mAd731_2 CB@4_mAd732_1 CB@4_mAd732_2 CB@4_mAd733_1 CB@4_mAd733_2 CB@4_mAd734_1 CB@4_mAd734_2 CB@4_mAd735_1 CB@4_mAd735_2 CB@4_mAd736_1 CB@4_mAd736_2 CB@4_mAd737_1 CB@4_mAd737_2 CB@4_mAd740_1 CB@4_mAd740_2 CB@4_mAd741_1 CB@4_mAd741_2 CB@4_mAd742_1 CB@4_mAd742_2 CB@4_mAd743_1 CB@4_mAd743_2 CB@4_mAd744_1 
+CB@4_mAd744_2 CB@4_mAd745_1 CB@4_mAd745_2 CB@4_mAd746_1 CB@4_mAd746_2 CB@4_mAd747_1 CB@4_mAd747_2 CB@4_mAd750_1 CB@4_mAd750_2 CB@4_mAd751_1 CB@4_mAd751_2 CB@4_mAd752_1 CB@4_mAd752_2 CB@4_mAd753_1 CB@4_mAd753_2 CB@4_mAd754_1 CB@4_mAd754_2 CB@4_mAd755_1 CB@4_mAd755_2 CB@4_mAd756_1 CB@4_mAd756_2 CB@4_mAd757_1 CB@4_mAd757_2 CB@4_mAd760_1 CB@4_mAd760_2 CB@4_mAd761_1 CB@4_mAd761_2 CB@4_mAd762_1 CB@4_mAd762_2 CB@4_mAd763_1 CB@4_mAd763_2 CB@4_mAd764_1 CB@4_mAd764_2 CB@4_mAd765_1 CB@4_mAd765_2 CB@4_mAd766_1 
+CB@4_mAd766_2 CB@4_mAd767_1 CB@4_mAd767_2 CB@4_mAd771_1 CB@4_mAd771_2 CB@4_mAd772_1 CB@4_mAd772_2 CB@4_mAd773_1 CB@4_mAd773_2 CB@4_mAd774_1 CB@4_mAd774_2 CB@4_mAd775_1 CB@4_mAd775_2 CB@4_mAd776_1 CB@4_mAd776_2 CB@4_mAd777_1 CB@4_mAd777_2 CB@4_X0 CB@4_X1 CB@4_X10 CB@4_X11 CB@4_X12 CB@4_X13 CB@4_X2 CB@4_X3 CB@4_X4 CB@4_X5 CB@4_X6 CB@4_X7 CB@4_X8 CB@4_X9 CB@4_Y1 CB@4_Y10 CB@4_Y11 CB@4_Y12 CB@4_Y2 CB@4_Y3 CB@4_Y4 CB@4_Y5 CB@4_Y6 CB@4_Y7 CB@4_Y8 CB@4_Y9 CB@4_Z1 CB@4_Z10 CB@4_Z11 CB@4_Z12 CB@4_Z2 CB@4_Z3 CB@4_Z4 
+CB@4_Z5 CB@4_Z6 CB@4_Z7 CB@4_Z8 CB@4_Z9 _5400TP094__CB
XCB@5 CB@5_K0 CB@5_K1 CB@5_K10 CB@5_K11 CB@5_K12 CB@5_K13 CB@5_K2 CB@5_K3 CB@5_K4 CB@5_K5 CB@5_K6 CB@5_K7 CB@5_K8 CB@5_K9 CB@5_mAd000_1 CB@5_mAd000_2 CB@5_mAd001_1 CB@5_mAd001_2 CB@5_mAd002_1 CB@5_mAd002_2 CB@5_mAd003_1 CB@5_mAd003_2 CB@5_mAd004_1 CB@5_mAd004_2 CB@5_mAd005_1 CB@5_mAd005_2 CB@5_mAd006_1 CB@5_mAd006_2 CB@5_mAd007_1 CB@5_mAd007_2 CB@5_mAd010_1 CB@5_mAd010_2 CB@5_mAd011_1 CB@5_mAd011_2 CB@5_mAd012_1 CB@5_mAd012_2 CB@5_mAd013_1 CB@5_mAd013_2 CB@5_mAd014_1 CB@5_mAd014_2 CB@5_mAd015_1 
+CB@5_mAd015_2 CB@5_mAd016_1 CB@5_mAd016_2 CB@5_mAd017_1 CB@5_mAd017_2 CB@5_mAd020_1 CB@5_mAd020_2 CB@5_mAd021_1 CB@5_mAd021_2 CB@5_mAd022_1 CB@5_mAd022_2 CB@5_mAd023_1 CB@5_mAd023_2 CB@5_mAd024_1 CB@5_mAd024_2 CB@5_mAd025_1 CB@5_mAd025_2 CB@5_mAd026_1 CB@5_mAd026_2 CB@5_mAd027_1 CB@5_mAd027_2 CB@5_mAd030_1 CB@5_mAd030_2 CB@5_mAd031_1 CB@5_mAd031_2 CB@5_mAd032_1 CB@5_mAd032_2 CB@5_mAd033_1 CB@5_mAd033_2 CB@5_mAd034_1 CB@5_mAd034_2 CB@5_mAd035_1 CB@5_mAd035_2 CB@5_mAd036_1 CB@5_mAd036_2 CB@5_mAd037_1 
+CB@5_mAd037_2 CB@5_mAd040_1 CB@5_mAd040_2 CB@5_mAd041_1 CB@5_mAd041_2 CB@5_mAd042_1 CB@5_mAd042_2 CB@5_mAd043_1 CB@5_mAd043_2 CB@5_mAd044_1 CB@5_mAd044_2 CB@5_mAd045_1 CB@5_mAd045_2 CB@5_mAd046_1 CB@5_mAd046_2 CB@5_mAd047_1 CB@5_mAd047_2 CB@5_mAd050_1 CB@5_mAd050_2 CB@5_mAd051_1 CB@5_mAd051_2 CB@5_mAd052_1 CB@5_mAd052_2 CB@5_mAd053_1 CB@5_mAd053_2 CB@5_mAd054_1 CB@5_mAd054_2 CB@5_mAd055_1 CB@5_mAd055_2 CB@5_mAd056_1 CB@5_mAd056_2 CB@5_mAd057_1 CB@5_mAd057_2 CB@5_mAd060_1 CB@5_mAd060_2 CB@5_mAd066_1 
+CB@5_mAd066_2 CB@5_mAd067_1 CB@5_mAd067_2 CB@5_mAd100_1 CB@5_mAd100_2 CB@5_mAd101_1 CB@5_mAd101_2 CB@5_mAd102_1 CB@5_mAd102_2 CB@5_mAd110_1 CB@5_mAd110_2 CB@5_mAd111_1 CB@5_mAd111_2 CB@5_mAd112_1 CB@5_mAd112_2 CB@5_mAd113_1 CB@5_mAd113_2 CB@5_mAd114_1 CB@5_mAd114_2 CB@5_mAd115_1 CB@5_mAd115_2 CB@5_mAd116_1 CB@5_mAd116_2 CB@5_mAd117_1 CB@5_mAd117_2 CB@5_mAd120_1 CB@5_mAd120_2 CB@5_mAd121_1 CB@5_mAd121_2 CB@5_mAd122_1 CB@5_mAd122_2 CB@5_mAd123_1 CB@5_mAd123_2 CB@5_mAd124_1 CB@5_mAd124_2 CB@5_mAd125_1 
+CB@5_mAd125_2 CB@5_mAd126_1 CB@5_mAd126_2 CB@5_mAd127_1 CB@5_mAd127_2 CB@5_mAd130_1 CB@5_mAd130_2 CB@5_mAd131_1 CB@5_mAd131_2 CB@5_mAd132_1 CB@5_mAd132_2 CB@5_mAd133_1 CB@5_mAd133_2 CB@5_mAd134_1 CB@5_mAd134_2 CB@5_mAd135_1 CB@5_mAd135_2 CB@5_mAd136_1 CB@5_mAd136_2 CB@5_mAd137_1 CB@5_mAd137_2 CB@5_mAd140_1 CB@5_mAd140_2 CB@5_mAd141_1 CB@5_mAd141_2 CB@5_mAd142_1 CB@5_mAd142_2 CB@5_mAd143_1 CB@5_mAd143_2 CB@5_mAd144_1 CB@5_mAd144_2 CB@5_mAd145_1 CB@5_mAd145_2 CB@5_mAd146_1 CB@5_mAd146_2 CB@5_mAd147_1 
+CB@5_mAd147_2 CB@5_mAd150_1 CB@5_mAd150_2 CB@5_mAd151_1 CB@5_mAd151_2 CB@5_mAd152_1 CB@5_mAd152_2 CB@5_mAd153_1 CB@5_mAd153_2 CB@5_mAd154_1 CB@5_mAd154_2 CB@5_mAd155_1 CB@5_mAd155_2 CB@5_mAd156_1 CB@5_mAd156_2 CB@5_mAd157_1 CB@5_mAd157_2 CB@5_mAd160_1 CB@5_mAd160_2 CB@5_mAd161_1 CB@5_mAd161_2 CB@5_mAd162_1 CB@5_mAd162_2 CB@5_mAd163_1 CB@5_mAd163_2 CB@5_mAd164_1 CB@5_mAd164_2 CB@5_mAd165_1 CB@5_mAd165_2 CB@5_mAd166_1 CB@5_mAd166_2 CB@5_mAd167_1 CB@5_mAd167_2 CB@5_mAd170_1 CB@5_mAd170_2 CB@5_mAd171_1 
+CB@5_mAd171_2 CB@5_mAd172_1 CB@5_mAd172_2 CB@5_mAd173_1 CB@5_mAd173_2 CB@5_mAd175_1 CB@5_mAd175_2 CB@5_mAd176_1 CB@5_mAd176_2 CB@5_mAd177_1 CB@5_mAd177_2 CB@5_mAd200_1 CB@5_mAd200_2 CB@5_mAd201_1 CB@5_mAd201_2 CB@5_mAd202_1 CB@5_mAd202_2 CB@5_mAd204_1 CB@5_mAd204_2 CB@5_mAd205_1 CB@5_mAd205_2 CB@5_mAd206_1 CB@5_mAd206_2 CB@5_mAd207_1 CB@5_mAd207_2 CB@5_mAd210_1 CB@5_mAd210_2 CB@5_mAd211_1 CB@5_mAd211_2 CB@5_mAd212_1 CB@5_mAd212_2 CB@5_mAd213_1 CB@5_mAd213_2 CB@5_mAd214_1 CB@5_mAd214_2 CB@5_mAd215_1 
+CB@5_mAd215_2 CB@5_mAd216_1 CB@5_mAd216_2 CB@5_mAd217_1 CB@5_mAd217_2 CB@5_mAd220_1 CB@5_mAd220_2 CB@5_mAd221_1 CB@5_mAd221_2 CB@5_mAd222_1 CB@5_mAd222_2 CB@5_mAd223_1 CB@5_mAd223_2 CB@5_mAd224_1 CB@5_mAd224_2 CB@5_mAd225_1 CB@5_mAd225_2 CB@5_mAd226_1 CB@5_mAd226_2 CB@5_mAd227_1 CB@5_mAd227_2 CB@5_mAd230_1 CB@5_mAd230_2 CB@5_mAd231_1 CB@5_mAd231_2 CB@5_mAd232_1 CB@5_mAd232_2 CB@5_mAd233_1 CB@5_mAd233_2 CB@5_mAd234_1 CB@5_mAd234_2 CB@5_mAd235_1 CB@5_mAd235_2 CB@5_mAd236_1 CB@5_mAd236_2 CB@5_mAd237_1 
+CB@5_mAd237_2 CB@5_mAd240_1 CB@5_mAd240_2 CB@5_mAd241_1 CB@5_mAd241_2 CB@5_mAd242_1 CB@5_mAd242_2 CB@5_mAd243_1 CB@5_mAd243_2 CB@5_mAd244_1 CB@5_mAd244_2 CB@5_mAd245_1 CB@5_mAd245_2 CB@5_mAd246_1 CB@5_mAd246_2 CB@5_mAd247_1 CB@5_mAd247_2 CB@5_mAd250_1 CB@5_mAd250_2 CB@5_mAd251_1 CB@5_mAd251_2 CB@5_mAd252_1 CB@5_mAd252_2 CB@5_mAd253_1 CB@5_mAd253_2 CB@5_mAd254_1 CB@5_mAd254_2 CB@5_mAd255_1 CB@5_mAd255_2 CB@5_mAd256_1 CB@5_mAd256_2 CB@5_mAd257_1 CB@5_mAd257_2 CB@5_mAd260_1 CB@5_mAd260_2 CB@5_mAd261_1 
+CB@5_mAd261_2 CB@5_mAd262_1 CB@5_mAd262_2 CB@5_mAd263_1 CB@5_mAd263_2 CB@5_mAd264_1 CB@5_mAd264_2 CB@5_mAd265_1 CB@5_mAd265_2 CB@5_mAd266_1 CB@5_mAd266_2 CB@5_mAd267_1 CB@5_mAd267_2 CB@5_mAd275_1 CB@5_mAd275_2 CB@5_mAd276_1 CB@5_mAd276_2 CB@5_mAd277_1 CB@5_mAd277_2 CB@5_mAd300_1 CB@5_mAd300_2 CB@5_mAd310_1 CB@5_mAd310_2 CB@5_mAd311_1 CB@5_mAd311_2 CB@5_mAd317_1 CB@5_mAd317_2 CB@5_mAd320_1 CB@5_mAd320_2 CB@5_mAd321_1 CB@5_mAd321_2 CB@5_mAd322_1 CB@5_mAd322_2 CB@5_mAd323_1 CB@5_mAd323_2 CB@5_mAd324_1 
+CB@5_mAd324_2 CB@5_mAd325_1 CB@5_mAd325_2 CB@5_mAd326_1 CB@5_mAd326_2 CB@5_mAd327_1 CB@5_mAd327_2 CB@5_mAd330_1 CB@5_mAd330_2 CB@5_mAd331_1 CB@5_mAd331_2 CB@5_mAd332_1 CB@5_mAd332_2 CB@5_mAd333_1 CB@5_mAd333_2 CB@5_mAd334_1 CB@5_mAd334_2 CB@5_mAd335_1 CB@5_mAd335_2 CB@5_mAd336_1 CB@5_mAd336_2 CB@5_mAd337_1 CB@5_mAd337_2 CB@5_mAd340_1 CB@5_mAd340_2 CB@5_mAd341_1 CB@5_mAd341_2 CB@5_mAd342_1 CB@5_mAd342_2 CB@5_mAd343_1 CB@5_mAd343_2 CB@5_mAd344_1 CB@5_mAd344_2 CB@5_mAd345_1 CB@5_mAd345_2 CB@5_mAd346_1 
+CB@5_mAd346_2 CB@5_mAd347_1 CB@5_mAd347_2 CB@5_mAd350_1 CB@5_mAd350_2 CB@5_mAd351_1 CB@5_mAd351_2 CB@5_mAd352_1 CB@5_mAd352_2 CB@5_mAd353_1 CB@5_mAd353_2 CB@5_mAd354_1 CB@5_mAd354_2 CB@5_mAd355_1 CB@5_mAd355_2 CB@5_mAd356_1 CB@5_mAd356_2 CB@5_mAd357_1 CB@5_mAd357_2 CB@5_mAd360_1 CB@5_mAd360_2 CB@5_mAd361_1 CB@5_mAd361_2 CB@5_mAd362_1 CB@5_mAd362_2 CB@5_mAd363_1 CB@5_mAd363_2 CB@5_mAd364_1 CB@5_mAd364_2 CB@5_mAd365_1 CB@5_mAd365_2 CB@5_mAd366_1 CB@5_mAd366_2 CB@5_mAd367_1 CB@5_mAd367_2 CB@5_mAd371_1 
+CB@5_mAd371_2 CB@5_mAd372_1 CB@5_mAd372_2 CB@5_mAd373_1 CB@5_mAd373_2 CB@5_mAd374_1 CB@5_mAd374_2 CB@5_mAd375_1 CB@5_mAd375_2 CB@5_mAd376_1 CB@5_mAd376_2 CB@5_mAd377_1 CB@5_mAd377_2 CB@5_mAd400_1 CB@5_mAd400_2 CB@5_mAd401_1 CB@5_mAd401_2 CB@5_mAd402_1 CB@5_mAd402_2 CB@5_mAd403_1 CB@5_mAd403_2 CB@5_mAd404_1 CB@5_mAd404_2 CB@5_mAd405_1 CB@5_mAd405_2 CB@5_mAd406_1 CB@5_mAd406_2 CB@5_mAd407_1 CB@5_mAd407_2 CB@5_mAd410_1 CB@5_mAd410_2 CB@5_mAd411_1 CB@5_mAd411_2 CB@5_mAd412_1 CB@5_mAd412_2 CB@5_mAd413_1 
+CB@5_mAd413_2 CB@5_mAd414_1 CB@5_mAd414_2 CB@5_mAd415_1 CB@5_mAd415_2 CB@5_mAd416_1 CB@5_mAd416_2 CB@5_mAd417_1 CB@5_mAd417_2 CB@5_mAd420_1 CB@5_mAd420_2 CB@5_mAd421_1 CB@5_mAd421_2 CB@5_mAd422_1 CB@5_mAd422_2 CB@5_mAd423_1 CB@5_mAd423_2 CB@5_mAd424_1 CB@5_mAd424_2 CB@5_mAd425_1 CB@5_mAd425_2 CB@5_mAd426_1 CB@5_mAd426_2 CB@5_mAd427_1 CB@5_mAd427_2 CB@5_mAd430_1 CB@5_mAd430_2 CB@5_mAd431_1 CB@5_mAd431_2 CB@5_mAd432_1 CB@5_mAd432_2 CB@5_mAd433_1 CB@5_mAd433_2 CB@5_mAd434_1 CB@5_mAd434_2 CB@5_mAd435_1 
+CB@5_mAd435_2 CB@5_mAd436_1 CB@5_mAd436_2 CB@5_mAd437_1 CB@5_mAd437_2 CB@5_mAd440_1 CB@5_mAd440_2 CB@5_mAd441_1 CB@5_mAd441_2 CB@5_mAd442_1 CB@5_mAd442_2 CB@5_mAd443_1 CB@5_mAd443_2 CB@5_mAd444_1 CB@5_mAd444_2 CB@5_mAd445_1 CB@5_mAd445_2 CB@5_mAd446_1 CB@5_mAd446_2 CB@5_mAd447_1 CB@5_mAd447_2 CB@5_mAd450_1 CB@5_mAd450_2 CB@5_mAd451_1 CB@5_mAd451_2 CB@5_mAd452_1 CB@5_mAd452_2 CB@5_mAd453_1 CB@5_mAd453_2 CB@5_mAd454_1 CB@5_mAd454_2 CB@5_mAd455_1 CB@5_mAd455_2 CB@5_mAd456_1 CB@5_mAd456_2 CB@5_mAd457_1 
+CB@5_mAd457_2 CB@5_mAd460_1 CB@5_mAd460_2 CB@5_mAd466_1 CB@5_mAd466_2 CB@5_mAd467_1 CB@5_mAd467_2 CB@5_mAd500_1 CB@5_mAd500_2 CB@5_mAd501_1 CB@5_mAd501_2 CB@5_mAd502_1 CB@5_mAd502_2 CB@5_mAd508_1 CB@5_mAd508_2 CB@5_mAd509_1 CB@5_mAd509_2 CB@5_mAd512_1 CB@5_mAd512_2 CB@5_mAd513_1 CB@5_mAd513_2 CB@5_mAd514_1 CB@5_mAd514_2 CB@5_mAd515_1 CB@5_mAd515_2 CB@5_mAd516_1 CB@5_mAd516_2 CB@5_mAd517_1 CB@5_mAd517_2 CB@5_mAd520_1 CB@5_mAd520_2 CB@5_mAd521_1 CB@5_mAd521_2 CB@5_mAd522_1 CB@5_mAd522_2 CB@5_mAd523_1 
+CB@5_mAd523_2 CB@5_mAd524_1 CB@5_mAd524_2 CB@5_mAd525_1 CB@5_mAd525_2 CB@5_mAd526_1 CB@5_mAd526_2 CB@5_mAd527_1 CB@5_mAd527_2 CB@5_mAd530_1 CB@5_mAd530_2 CB@5_mAd531_1 CB@5_mAd531_2 CB@5_mAd532_1 CB@5_mAd532_2 CB@5_mAd533_1 CB@5_mAd533_2 CB@5_mAd534_1 CB@5_mAd534_2 CB@5_mAd535_1 CB@5_mAd535_2 CB@5_mAd536_1 CB@5_mAd536_2 CB@5_mAd537_1 CB@5_mAd537_2 CB@5_mAd540_1 CB@5_mAd540_2 CB@5_mAd541_1 CB@5_mAd541_2 CB@5_mAd542_1 CB@5_mAd542_2 CB@5_mAd543_1 CB@5_mAd543_2 CB@5_mAd544_1 CB@5_mAd544_2 CB@5_mAd545_1 
+CB@5_mAd545_2 CB@5_mAd546_1 CB@5_mAd546_2 CB@5_mAd547_1 CB@5_mAd547_2 CB@5_mAd550_1 CB@5_mAd550_2 CB@5_mAd551_1 CB@5_mAd551_2 CB@5_mAd552_1 CB@5_mAd552_2 CB@5_mAd553_1 CB@5_mAd553_2 CB@5_mAd554_1 CB@5_mAd554_2 CB@5_mAd555_1 CB@5_mAd555_2 CB@5_mAd556_1 CB@5_mAd556_2 CB@5_mAd557_1 CB@5_mAd557_2 CB@5_mAd560_1 CB@5_mAd560_2 CB@5_mAd561_1 CB@5_mAd561_2 CB@5_mAd562_1 CB@5_mAd562_2 CB@5_mAd563_1 CB@5_mAd563_2 CB@5_mAd564_1 CB@5_mAd564_2 CB@5_mAd565_1 CB@5_mAd565_2 CB@5_mAd566_1 CB@5_mAd566_2 CB@5_mAd567_1 
+CB@5_mAd567_2 CB@5_mAd570_1 CB@5_mAd570_2 CB@5_mAd571_1 CB@5_mAd571_2 CB@5_mAd572_1 CB@5_mAd572_2 CB@5_mAd573_1 CB@5_mAd573_2 CB@5_mAd575_1 CB@5_mAd575_2 CB@5_mAd576_1 CB@5_mAd576_2 CB@5_mAd577_1 CB@5_mAd577_2 CB@5_mAd600_1 CB@5_mAd600_2 CB@5_mAd601_1 CB@5_mAd601_2 CB@5_mAd602_1 CB@5_mAd602_2 CB@5_mAd604_1 CB@5_mAd604_2 CB@5_mAd605_1 CB@5_mAd605_2 CB@5_mAd606_1 CB@5_mAd606_2 CB@5_mAd607_1 CB@5_mAd607_2 CB@5_mAd610_1 CB@5_mAd610_2 CB@5_mAd611_1 CB@5_mAd611_2 CB@5_mAd612_1 CB@5_mAd612_2 CB@5_mAd613_1 
+CB@5_mAd613_2 CB@5_mAd614_1 CB@5_mAd614_2 CB@5_mAd615_1 CB@5_mAd615_2 CB@5_mAd616_1 CB@5_mAd616_2 CB@5_mAd617_1 CB@5_mAd617_2 CB@5_mAd620_1 CB@5_mAd620_2 CB@5_mAd621_1 CB@5_mAd621_2 CB@5_mAd622_1 CB@5_mAd622_2 CB@5_mAd623_1 CB@5_mAd623_2 CB@5_mAd624_1 CB@5_mAd624_2 CB@5_mAd625_1 CB@5_mAd625_2 CB@5_mAd626_1 CB@5_mAd626_2 CB@5_mAd627_1 CB@5_mAd627_2 CB@5_mAd630_1 CB@5_mAd630_2 CB@5_mAd631_1 CB@5_mAd631_2 CB@5_mAd632_1 CB@5_mAd632_2 CB@5_mAd633_1 CB@5_mAd633_2 CB@5_mAd634_1 CB@5_mAd634_2 CB@5_mAd635_1 
+CB@5_mAd635_2 CB@5_mAd636_1 CB@5_mAd636_2 CB@5_mAd637_1 CB@5_mAd637_2 CB@5_mAd640_1 CB@5_mAd640_2 CB@5_mAd641_1 CB@5_mAd641_2 CB@5_mAd642_1 CB@5_mAd642_2 CB@5_mAd643_1 CB@5_mAd643_2 CB@5_mAd644_1 CB@5_mAd644_2 CB@5_mAd645_1 CB@5_mAd645_2 CB@5_mAd646_1 CB@5_mAd646_2 CB@5_mAd647_1 CB@5_mAd647_2 CB@5_mAd650_1 CB@5_mAd650_2 CB@5_mAd651_1 CB@5_mAd651_2 CB@5_mAd652_1 CB@5_mAd652_2 CB@5_mAd653_1 CB@5_mAd653_2 CB@5_mAd654_1 CB@5_mAd654_2 CB@5_mAd655_1 CB@5_mAd655_2 CB@5_mAd656_1 CB@5_mAd656_2 CB@5_mAd657_1 
+CB@5_mAd657_2 CB@5_mAd660_1 CB@5_mAd660_2 CB@5_mAd661_1 CB@5_mAd661_2 CB@5_mAd662_1 CB@5_mAd662_2 CB@5_mAd663_1 CB@5_mAd663_2 CB@5_mAd664_1 CB@5_mAd664_2 CB@5_mAd665_1 CB@5_mAd665_2 CB@5_mAd666_1 CB@5_mAd666_2 CB@5_mAd667_1 CB@5_mAd667_2 CB@5_mAd675_1 CB@5_mAd675_2 CB@5_mAd676_1 CB@5_mAd676_2 CB@5_mAd677_1 CB@5_mAd677_2 CB@5_mAd700_1 CB@5_mAd700_2 CB@5_mAd710_1 CB@5_mAd710_2 CB@5_mAd711_1 CB@5_mAd711_2 CB@5_mAd717_1 CB@5_mAd717_2 CB@5_mAd720_1 CB@5_mAd720_2 CB@5_mAd721_1 CB@5_mAd721_2 CB@5_mAd722_1 
+CB@5_mAd722_2 CB@5_mAd723_1 CB@5_mAd723_2 CB@5_mAd724_1 CB@5_mAd724_2 CB@5_mAd725_1 CB@5_mAd725_2 CB@5_mAd726_1 CB@5_mAd726_2 CB@5_mAd727_1 CB@5_mAd727_2 CB@5_mAd730_1 CB@5_mAd730_2 CB@5_mAd731_1 CB@5_mAd731_2 CB@5_mAd732_1 CB@5_mAd732_2 CB@5_mAd733_1 CB@5_mAd733_2 CB@5_mAd734_1 CB@5_mAd734_2 CB@5_mAd735_1 CB@5_mAd735_2 CB@5_mAd736_1 CB@5_mAd736_2 CB@5_mAd737_1 CB@5_mAd737_2 CB@5_mAd740_1 CB@5_mAd740_2 CB@5_mAd741_1 CB@5_mAd741_2 CB@5_mAd742_1 CB@5_mAd742_2 CB@5_mAd743_1 CB@5_mAd743_2 CB@5_mAd744_1 
+CB@5_mAd744_2 CB@5_mAd745_1 CB@5_mAd745_2 CB@5_mAd746_1 CB@5_mAd746_2 CB@5_mAd747_1 CB@5_mAd747_2 CB@5_mAd750_1 CB@5_mAd750_2 CB@5_mAd751_1 CB@5_mAd751_2 CB@5_mAd752_1 CB@5_mAd752_2 CB@5_mAd753_1 CB@5_mAd753_2 CB@5_mAd754_1 CB@5_mAd754_2 CB@5_mAd755_1 CB@5_mAd755_2 CB@5_mAd756_1 CB@5_mAd756_2 CB@5_mAd757_1 CB@5_mAd757_2 CB@5_mAd760_1 CB@5_mAd760_2 CB@5_mAd761_1 CB@5_mAd761_2 CB@5_mAd762_1 CB@5_mAd762_2 CB@5_mAd763_1 CB@5_mAd763_2 CB@5_mAd764_1 CB@5_mAd764_2 CB@5_mAd765_1 CB@5_mAd765_2 CB@5_mAd766_1 
+CB@5_mAd766_2 CB@5_mAd767_1 CB@5_mAd767_2 CB@5_mAd771_1 CB@5_mAd771_2 CB@5_mAd772_1 CB@5_mAd772_2 CB@5_mAd773_1 CB@5_mAd773_2 CB@5_mAd774_1 CB@5_mAd774_2 CB@5_mAd775_1 CB@5_mAd775_2 CB@5_mAd776_1 CB@5_mAd776_2 CB@5_mAd777_1 CB@5_mAd777_2 CB@5_X0 CB@5_X1 CB@5_X10 CB@5_X11 CB@5_X12 CB@5_X13 CB@5_X2 CB@5_X3 CB@5_X4 CB@5_X5 CB@5_X6 CB@5_X7 CB@5_X8 CB@5_X9 CB@5_Y1 CB@5_Y10 CB@5_Y11 CB@5_Y12 CB@5_Y2 CB@5_Y3 CB@5_Y4 CB@5_Y5 CB@5_Y6 CB@5_Y7 CB@5_Y8 CB@5_Y9 CB@5_Z1 CB@5_Z10 CB@5_Z11 CB@5_Z12 CB@5_Z2 CB@5_Z3 CB@5_Z4 
+CB@5_Z5 CB@5_Z6 CB@5_Z7 CB@5_Z8 CB@5_Z9 _5400TP094__CB
XCB@6 CB@6_K0 CB@6_K1 CB@6_K10 CB@6_K11 CB@6_K12 CB@6_K13 CB@6_K2 CB@6_K3 CB@6_K4 CB@6_K5 CB@6_K6 CB@6_K7 CB@6_K8 CB@6_K9 CB@6_mAd000_1 CB@6_mAd000_2 CB@6_mAd001_1 CB@6_mAd001_2 CB@6_mAd002_1 CB@6_mAd002_2 CB@6_mAd003_1 CB@6_mAd003_2 CB@6_mAd004_1 CB@6_mAd004_2 CB@6_mAd005_1 CB@6_mAd005_2 CB@6_mAd006_1 CB@6_mAd006_2 CB@6_mAd007_1 CB@6_mAd007_2 CB@6_mAd010_1 CB@6_mAd010_2 CB@6_mAd011_1 CB@6_mAd011_2 CB@6_mAd012_1 CB@6_mAd012_2 CB@6_mAd013_1 CB@6_mAd013_2 CB@6_mAd014_1 CB@6_mAd014_2 CB@6_mAd015_1 
+CB@6_mAd015_2 CB@6_mAd016_1 CB@6_mAd016_2 CB@6_mAd017_1 CB@6_mAd017_2 CB@6_mAd020_1 CB@6_mAd020_2 CB@6_mAd021_1 CB@6_mAd021_2 CB@6_mAd022_1 CB@6_mAd022_2 CB@6_mAd023_1 CB@6_mAd023_2 CB@6_mAd024_1 CB@6_mAd024_2 CB@6_mAd025_1 CB@6_mAd025_2 CB@6_mAd026_1 CB@6_mAd026_2 CB@6_mAd027_1 CB@6_mAd027_2 CB@6_mAd030_1 CB@6_mAd030_2 CB@6_mAd031_1 CB@6_mAd031_2 CB@6_mAd032_1 CB@6_mAd032_2 CB@6_mAd033_1 CB@6_mAd033_2 CB@6_mAd034_1 CB@6_mAd034_2 CB@6_mAd035_1 CB@6_mAd035_2 CB@6_mAd036_1 CB@6_mAd036_2 CB@6_mAd037_1 
+CB@6_mAd037_2 CB@6_mAd040_1 CB@6_mAd040_2 CB@6_mAd041_1 CB@6_mAd041_2 CB@6_mAd042_1 CB@6_mAd042_2 CB@6_mAd043_1 CB@6_mAd043_2 CB@6_mAd044_1 CB@6_mAd044_2 CB@6_mAd045_1 CB@6_mAd045_2 CB@6_mAd046_1 CB@6_mAd046_2 CB@6_mAd047_1 CB@6_mAd047_2 CB@6_mAd050_1 CB@6_mAd050_2 CB@6_mAd051_1 CB@6_mAd051_2 CB@6_mAd052_1 CB@6_mAd052_2 CB@6_mAd053_1 CB@6_mAd053_2 CB@6_mAd054_1 CB@6_mAd054_2 CB@6_mAd055_1 CB@6_mAd055_2 CB@6_mAd056_1 CB@6_mAd056_2 CB@6_mAd057_1 CB@6_mAd057_2 CB@6_mAd060_1 CB@6_mAd060_2 CB@6_mAd066_1 
+CB@6_mAd066_2 CB@6_mAd067_1 CB@6_mAd067_2 CB@6_mAd100_1 CB@6_mAd100_2 CB@6_mAd101_1 CB@6_mAd101_2 CB@6_mAd102_1 CB@6_mAd102_2 CB@6_mAd110_1 CB@6_mAd110_2 CB@6_mAd111_1 CB@6_mAd111_2 CB@6_mAd112_1 CB@6_mAd112_2 CB@6_mAd113_1 CB@6_mAd113_2 CB@6_mAd114_1 CB@6_mAd114_2 CB@6_mAd115_1 CB@6_mAd115_2 CB@6_mAd116_1 CB@6_mAd116_2 CB@6_mAd117_1 CB@6_mAd117_2 CB@6_mAd120_1 CB@6_mAd120_2 CB@6_mAd121_1 CB@6_mAd121_2 CB@6_mAd122_1 CB@6_mAd122_2 CB@6_mAd123_1 CB@6_mAd123_2 CB@6_mAd124_1 CB@6_mAd124_2 CB@6_mAd125_1 
+CB@6_mAd125_2 CB@6_mAd126_1 CB@6_mAd126_2 CB@6_mAd127_1 CB@6_mAd127_2 CB@6_mAd130_1 CB@6_mAd130_2 CB@6_mAd131_1 CB@6_mAd131_2 CB@6_mAd132_1 CB@6_mAd132_2 CB@6_mAd133_1 CB@6_mAd133_2 CB@6_mAd134_1 CB@6_mAd134_2 CB@6_mAd135_1 CB@6_mAd135_2 CB@6_mAd136_1 CB@6_mAd136_2 CB@6_mAd137_1 CB@6_mAd137_2 CB@6_mAd140_1 CB@6_mAd140_2 CB@6_mAd141_1 CB@6_mAd141_2 CB@6_mAd142_1 CB@6_mAd142_2 CB@6_mAd143_1 CB@6_mAd143_2 CB@6_mAd144_1 CB@6_mAd144_2 CB@6_mAd145_1 CB@6_mAd145_2 CB@6_mAd146_1 CB@6_mAd146_2 CB@6_mAd147_1 
+CB@6_mAd147_2 CB@6_mAd150_1 CB@6_mAd150_2 CB@6_mAd151_1 CB@6_mAd151_2 CB@6_mAd152_1 CB@6_mAd152_2 CB@6_mAd153_1 CB@6_mAd153_2 CB@6_mAd154_1 CB@6_mAd154_2 CB@6_mAd155_1 CB@6_mAd155_2 CB@6_mAd156_1 CB@6_mAd156_2 CB@6_mAd157_1 CB@6_mAd157_2 CB@6_mAd160_1 CB@6_mAd160_2 CB@6_mAd161_1 CB@6_mAd161_2 CB@6_mAd162_1 CB@6_mAd162_2 CB@6_mAd163_1 CB@6_mAd163_2 CB@6_mAd164_1 CB@6_mAd164_2 CB@6_mAd165_1 CB@6_mAd165_2 CB@6_mAd166_1 CB@6_mAd166_2 CB@6_mAd167_1 CB@6_mAd167_2 CB@6_mAd170_1 CB@6_mAd170_2 CB@6_mAd171_1 
+CB@6_mAd171_2 CB@6_mAd172_1 CB@6_mAd172_2 CB@6_mAd173_1 CB@6_mAd173_2 CB@6_mAd175_1 CB@6_mAd175_2 CB@6_mAd176_1 CB@6_mAd176_2 CB@6_mAd177_1 CB@6_mAd177_2 CB@6_mAd200_1 CB@6_mAd200_2 CB@6_mAd201_1 CB@6_mAd201_2 CB@6_mAd202_1 CB@6_mAd202_2 CB@6_mAd204_1 CB@6_mAd204_2 CB@6_mAd205_1 CB@6_mAd205_2 CB@6_mAd206_1 CB@6_mAd206_2 CB@6_mAd207_1 CB@6_mAd207_2 CB@6_mAd210_1 CB@6_mAd210_2 CB@6_mAd211_1 CB@6_mAd211_2 CB@6_mAd212_1 CB@6_mAd212_2 CB@6_mAd213_1 CB@6_mAd213_2 CB@6_mAd214_1 CB@6_mAd214_2 CB@6_mAd215_1 
+CB@6_mAd215_2 CB@6_mAd216_1 CB@6_mAd216_2 CB@6_mAd217_1 CB@6_mAd217_2 CB@6_mAd220_1 CB@6_mAd220_2 CB@6_mAd221_1 CB@6_mAd221_2 CB@6_mAd222_1 CB@6_mAd222_2 CB@6_mAd223_1 CB@6_mAd223_2 CB@6_mAd224_1 CB@6_mAd224_2 CB@6_mAd225_1 CB@6_mAd225_2 CB@6_mAd226_1 CB@6_mAd226_2 CB@6_mAd227_1 CB@6_mAd227_2 CB@6_mAd230_1 CB@6_mAd230_2 CB@6_mAd231_1 CB@6_mAd231_2 CB@6_mAd232_1 CB@6_mAd232_2 CB@6_mAd233_1 CB@6_mAd233_2 CB@6_mAd234_1 CB@6_mAd234_2 CB@6_mAd235_1 CB@6_mAd235_2 CB@6_mAd236_1 CB@6_mAd236_2 CB@6_mAd237_1 
+CB@6_mAd237_2 CB@6_mAd240_1 CB@6_mAd240_2 CB@6_mAd241_1 CB@6_mAd241_2 CB@6_mAd242_1 CB@6_mAd242_2 CB@6_mAd243_1 CB@6_mAd243_2 CB@6_mAd244_1 CB@6_mAd244_2 CB@6_mAd245_1 CB@6_mAd245_2 CB@6_mAd246_1 CB@6_mAd246_2 CB@6_mAd247_1 CB@6_mAd247_2 CB@6_mAd250_1 CB@6_mAd250_2 CB@6_mAd251_1 CB@6_mAd251_2 CB@6_mAd252_1 CB@6_mAd252_2 CB@6_mAd253_1 CB@6_mAd253_2 CB@6_mAd254_1 CB@6_mAd254_2 CB@6_mAd255_1 CB@6_mAd255_2 CB@6_mAd256_1 CB@6_mAd256_2 CB@6_mAd257_1 CB@6_mAd257_2 CB@6_mAd260_1 CB@6_mAd260_2 CB@6_mAd261_1 
+CB@6_mAd261_2 CB@6_mAd262_1 CB@6_mAd262_2 CB@6_mAd263_1 CB@6_mAd263_2 CB@6_mAd264_1 CB@6_mAd264_2 CB@6_mAd265_1 CB@6_mAd265_2 CB@6_mAd266_1 CB@6_mAd266_2 CB@6_mAd267_1 CB@6_mAd267_2 CB@6_mAd275_1 CB@6_mAd275_2 CB@6_mAd276_1 CB@6_mAd276_2 CB@6_mAd277_1 CB@6_mAd277_2 CB@6_mAd300_1 CB@6_mAd300_2 CB@6_mAd310_1 CB@6_mAd310_2 CB@6_mAd311_1 CB@6_mAd311_2 CB@6_mAd317_1 CB@6_mAd317_2 CB@6_mAd320_1 CB@6_mAd320_2 CB@6_mAd321_1 CB@6_mAd321_2 CB@6_mAd322_1 CB@6_mAd322_2 CB@6_mAd323_1 CB@6_mAd323_2 CB@6_mAd324_1 
+CB@6_mAd324_2 CB@6_mAd325_1 CB@6_mAd325_2 CB@6_mAd326_1 CB@6_mAd326_2 CB@6_mAd327_1 CB@6_mAd327_2 CB@6_mAd330_1 CB@6_mAd330_2 CB@6_mAd331_1 CB@6_mAd331_2 CB@6_mAd332_1 CB@6_mAd332_2 CB@6_mAd333_1 CB@6_mAd333_2 CB@6_mAd334_1 CB@6_mAd334_2 CB@6_mAd335_1 CB@6_mAd335_2 CB@6_mAd336_1 CB@6_mAd336_2 CB@6_mAd337_1 CB@6_mAd337_2 CB@6_mAd340_1 CB@6_mAd340_2 CB@6_mAd341_1 CB@6_mAd341_2 CB@6_mAd342_1 CB@6_mAd342_2 CB@6_mAd343_1 CB@6_mAd343_2 CB@6_mAd344_1 CB@6_mAd344_2 CB@6_mAd345_1 CB@6_mAd345_2 CB@6_mAd346_1 
+CB@6_mAd346_2 CB@6_mAd347_1 CB@6_mAd347_2 CB@6_mAd350_1 CB@6_mAd350_2 CB@6_mAd351_1 CB@6_mAd351_2 CB@6_mAd352_1 CB@6_mAd352_2 CB@6_mAd353_1 CB@6_mAd353_2 CB@6_mAd354_1 CB@6_mAd354_2 CB@6_mAd355_1 CB@6_mAd355_2 CB@6_mAd356_1 CB@6_mAd356_2 CB@6_mAd357_1 CB@6_mAd357_2 CB@6_mAd360_1 CB@6_mAd360_2 CB@6_mAd361_1 CB@6_mAd361_2 CB@6_mAd362_1 CB@6_mAd362_2 CB@6_mAd363_1 CB@6_mAd363_2 CB@6_mAd364_1 CB@6_mAd364_2 CB@6_mAd365_1 CB@6_mAd365_2 CB@6_mAd366_1 CB@6_mAd366_2 CB@6_mAd367_1 CB@6_mAd367_2 CB@6_mAd371_1 
+CB@6_mAd371_2 CB@6_mAd372_1 CB@6_mAd372_2 CB@6_mAd373_1 CB@6_mAd373_2 CB@6_mAd374_1 CB@6_mAd374_2 CB@6_mAd375_1 CB@6_mAd375_2 CB@6_mAd376_1 CB@6_mAd376_2 CB@6_mAd377_1 CB@6_mAd377_2 CB@6_mAd400_1 CB@6_mAd400_2 CB@6_mAd401_1 CB@6_mAd401_2 CB@6_mAd402_1 CB@6_mAd402_2 CB@6_mAd403_1 CB@6_mAd403_2 CB@6_mAd404_1 CB@6_mAd404_2 CB@6_mAd405_1 CB@6_mAd405_2 CB@6_mAd406_1 CB@6_mAd406_2 CB@6_mAd407_1 CB@6_mAd407_2 CB@6_mAd410_1 CB@6_mAd410_2 CB@6_mAd411_1 CB@6_mAd411_2 CB@6_mAd412_1 CB@6_mAd412_2 CB@6_mAd413_1 
+CB@6_mAd413_2 CB@6_mAd414_1 CB@6_mAd414_2 CB@6_mAd415_1 CB@6_mAd415_2 CB@6_mAd416_1 CB@6_mAd416_2 CB@6_mAd417_1 CB@6_mAd417_2 CB@6_mAd420_1 CB@6_mAd420_2 CB@6_mAd421_1 CB@6_mAd421_2 CB@6_mAd422_1 CB@6_mAd422_2 CB@6_mAd423_1 CB@6_mAd423_2 CB@6_mAd424_1 CB@6_mAd424_2 CB@6_mAd425_1 CB@6_mAd425_2 CB@6_mAd426_1 CB@6_mAd426_2 CB@6_mAd427_1 CB@6_mAd427_2 CB@6_mAd430_1 CB@6_mAd430_2 CB@6_mAd431_1 CB@6_mAd431_2 CB@6_mAd432_1 CB@6_mAd432_2 CB@6_mAd433_1 CB@6_mAd433_2 CB@6_mAd434_1 CB@6_mAd434_2 CB@6_mAd435_1 
+CB@6_mAd435_2 CB@6_mAd436_1 CB@6_mAd436_2 CB@6_mAd437_1 CB@6_mAd437_2 CB@6_mAd440_1 CB@6_mAd440_2 CB@6_mAd441_1 CB@6_mAd441_2 CB@6_mAd442_1 CB@6_mAd442_2 CB@6_mAd443_1 CB@6_mAd443_2 CB@6_mAd444_1 CB@6_mAd444_2 CB@6_mAd445_1 CB@6_mAd445_2 CB@6_mAd446_1 CB@6_mAd446_2 CB@6_mAd447_1 CB@6_mAd447_2 CB@6_mAd450_1 CB@6_mAd450_2 CB@6_mAd451_1 CB@6_mAd451_2 CB@6_mAd452_1 CB@6_mAd452_2 CB@6_mAd453_1 CB@6_mAd453_2 CB@6_mAd454_1 CB@6_mAd454_2 CB@6_mAd455_1 CB@6_mAd455_2 CB@6_mAd456_1 CB@6_mAd456_2 CB@6_mAd457_1 
+CB@6_mAd457_2 CB@6_mAd460_1 CB@6_mAd460_2 CB@6_mAd466_1 CB@6_mAd466_2 CB@6_mAd467_1 CB@6_mAd467_2 CB@6_mAd500_1 CB@6_mAd500_2 CB@6_mAd501_1 CB@6_mAd501_2 CB@6_mAd502_1 CB@6_mAd502_2 CB@6_mAd508_1 CB@6_mAd508_2 CB@6_mAd509_1 CB@6_mAd509_2 CB@6_mAd512_1 CB@6_mAd512_2 CB@6_mAd513_1 CB@6_mAd513_2 CB@6_mAd514_1 CB@6_mAd514_2 CB@6_mAd515_1 CB@6_mAd515_2 CB@6_mAd516_1 CB@6_mAd516_2 CB@6_mAd517_1 CB@6_mAd517_2 CB@6_mAd520_1 CB@6_mAd520_2 CB@6_mAd521_1 CB@6_mAd521_2 CB@6_mAd522_1 CB@6_mAd522_2 CB@6_mAd523_1 
+CB@6_mAd523_2 CB@6_mAd524_1 CB@6_mAd524_2 CB@6_mAd525_1 CB@6_mAd525_2 CB@6_mAd526_1 CB@6_mAd526_2 CB@6_mAd527_1 CB@6_mAd527_2 CB@6_mAd530_1 CB@6_mAd530_2 CB@6_mAd531_1 CB@6_mAd531_2 CB@6_mAd532_1 CB@6_mAd532_2 CB@6_mAd533_1 CB@6_mAd533_2 CB@6_mAd534_1 CB@6_mAd534_2 CB@6_mAd535_1 CB@6_mAd535_2 CB@6_mAd536_1 CB@6_mAd536_2 CB@6_mAd537_1 CB@6_mAd537_2 CB@6_mAd540_1 CB@6_mAd540_2 CB@6_mAd541_1 CB@6_mAd541_2 CB@6_mAd542_1 CB@6_mAd542_2 CB@6_mAd543_1 CB@6_mAd543_2 CB@6_mAd544_1 CB@6_mAd544_2 CB@6_mAd545_1 
+CB@6_mAd545_2 CB@6_mAd546_1 CB@6_mAd546_2 CB@6_mAd547_1 CB@6_mAd547_2 CB@6_mAd550_1 CB@6_mAd550_2 CB@6_mAd551_1 CB@6_mAd551_2 CB@6_mAd552_1 CB@6_mAd552_2 CB@6_mAd553_1 CB@6_mAd553_2 CB@6_mAd554_1 CB@6_mAd554_2 CB@6_mAd555_1 CB@6_mAd555_2 CB@6_mAd556_1 CB@6_mAd556_2 CB@6_mAd557_1 CB@6_mAd557_2 CB@6_mAd560_1 CB@6_mAd560_2 CB@6_mAd561_1 CB@6_mAd561_2 CB@6_mAd562_1 CB@6_mAd562_2 CB@6_mAd563_1 CB@6_mAd563_2 CB@6_mAd564_1 CB@6_mAd564_2 CB@6_mAd565_1 CB@6_mAd565_2 CB@6_mAd566_1 CB@6_mAd566_2 CB@6_mAd567_1 
+CB@6_mAd567_2 CB@6_mAd570_1 CB@6_mAd570_2 CB@6_mAd571_1 CB@6_mAd571_2 CB@6_mAd572_1 CB@6_mAd572_2 CB@6_mAd573_1 CB@6_mAd573_2 CB@6_mAd575_1 CB@6_mAd575_2 CB@6_mAd576_1 CB@6_mAd576_2 CB@6_mAd577_1 CB@6_mAd577_2 CB@6_mAd600_1 CB@6_mAd600_2 CB@6_mAd601_1 CB@6_mAd601_2 CB@6_mAd602_1 CB@6_mAd602_2 CB@6_mAd604_1 CB@6_mAd604_2 CB@6_mAd605_1 CB@6_mAd605_2 CB@6_mAd606_1 CB@6_mAd606_2 CB@6_mAd607_1 CB@6_mAd607_2 CB@6_mAd610_1 CB@6_mAd610_2 CB@6_mAd611_1 CB@6_mAd611_2 CB@6_mAd612_1 CB@6_mAd612_2 CB@6_mAd613_1 
+CB@6_mAd613_2 CB@6_mAd614_1 CB@6_mAd614_2 CB@6_mAd615_1 CB@6_mAd615_2 CB@6_mAd616_1 CB@6_mAd616_2 CB@6_mAd617_1 CB@6_mAd617_2 CB@6_mAd620_1 CB@6_mAd620_2 CB@6_mAd621_1 CB@6_mAd621_2 CB@6_mAd622_1 CB@6_mAd622_2 CB@6_mAd623_1 CB@6_mAd623_2 CB@6_mAd624_1 CB@6_mAd624_2 CB@6_mAd625_1 CB@6_mAd625_2 CB@6_mAd626_1 CB@6_mAd626_2 CB@6_mAd627_1 CB@6_mAd627_2 CB@6_mAd630_1 CB@6_mAd630_2 CB@6_mAd631_1 CB@6_mAd631_2 CB@6_mAd632_1 CB@6_mAd632_2 CB@6_mAd633_1 CB@6_mAd633_2 CB@6_mAd634_1 CB@6_mAd634_2 CB@6_mAd635_1 
+CB@6_mAd635_2 CB@6_mAd636_1 CB@6_mAd636_2 CB@6_mAd637_1 CB@6_mAd637_2 CB@6_mAd640_1 CB@6_mAd640_2 CB@6_mAd641_1 CB@6_mAd641_2 CB@6_mAd642_1 CB@6_mAd642_2 CB@6_mAd643_1 CB@6_mAd643_2 CB@6_mAd644_1 CB@6_mAd644_2 CB@6_mAd645_1 CB@6_mAd645_2 CB@6_mAd646_1 CB@6_mAd646_2 CB@6_mAd647_1 CB@6_mAd647_2 CB@6_mAd650_1 CB@6_mAd650_2 CB@6_mAd651_1 CB@6_mAd651_2 CB@6_mAd652_1 CB@6_mAd652_2 CB@6_mAd653_1 CB@6_mAd653_2 CB@6_mAd654_1 CB@6_mAd654_2 CB@6_mAd655_1 CB@6_mAd655_2 CB@6_mAd656_1 CB@6_mAd656_2 CB@6_mAd657_1 
+CB@6_mAd657_2 CB@6_mAd660_1 CB@6_mAd660_2 CB@6_mAd661_1 CB@6_mAd661_2 CB@6_mAd662_1 CB@6_mAd662_2 CB@6_mAd663_1 CB@6_mAd663_2 CB@6_mAd664_1 CB@6_mAd664_2 CB@6_mAd665_1 CB@6_mAd665_2 CB@6_mAd666_1 CB@6_mAd666_2 CB@6_mAd667_1 CB@6_mAd667_2 CB@6_mAd675_1 CB@6_mAd675_2 CB@6_mAd676_1 CB@6_mAd676_2 CB@6_mAd677_1 CB@6_mAd677_2 CB@6_mAd700_1 CB@6_mAd700_2 CB@6_mAd710_1 CB@6_mAd710_2 CB@6_mAd711_1 CB@6_mAd711_2 CB@6_mAd717_1 CB@6_mAd717_2 CB@6_mAd720_1 CB@6_mAd720_2 CB@6_mAd721_1 CB@6_mAd721_2 CB@6_mAd722_1 
+CB@6_mAd722_2 CB@6_mAd723_1 CB@6_mAd723_2 CB@6_mAd724_1 CB@6_mAd724_2 CB@6_mAd725_1 CB@6_mAd725_2 CB@6_mAd726_1 CB@6_mAd726_2 CB@6_mAd727_1 CB@6_mAd727_2 CB@6_mAd730_1 CB@6_mAd730_2 CB@6_mAd731_1 CB@6_mAd731_2 CB@6_mAd732_1 CB@6_mAd732_2 CB@6_mAd733_1 CB@6_mAd733_2 CB@6_mAd734_1 CB@6_mAd734_2 CB@6_mAd735_1 CB@6_mAd735_2 CB@6_mAd736_1 CB@6_mAd736_2 CB@6_mAd737_1 CB@6_mAd737_2 CB@6_mAd740_1 CB@6_mAd740_2 CB@6_mAd741_1 CB@6_mAd741_2 CB@6_mAd742_1 CB@6_mAd742_2 CB@6_mAd743_1 CB@6_mAd743_2 CB@6_mAd744_1 
+CB@6_mAd744_2 CB@6_mAd745_1 CB@6_mAd745_2 CB@6_mAd746_1 CB@6_mAd746_2 CB@6_mAd747_1 CB@6_mAd747_2 CB@6_mAd750_1 CB@6_mAd750_2 CB@6_mAd751_1 CB@6_mAd751_2 CB@6_mAd752_1 CB@6_mAd752_2 CB@6_mAd753_1 CB@6_mAd753_2 CB@6_mAd754_1 CB@6_mAd754_2 CB@6_mAd755_1 CB@6_mAd755_2 CB@6_mAd756_1 CB@6_mAd756_2 CB@6_mAd757_1 CB@6_mAd757_2 CB@6_mAd760_1 CB@6_mAd760_2 CB@6_mAd761_1 CB@6_mAd761_2 CB@6_mAd762_1 CB@6_mAd762_2 CB@6_mAd763_1 CB@6_mAd763_2 CB@6_mAd764_1 CB@6_mAd764_2 CB@6_mAd765_1 CB@6_mAd765_2 CB@6_mAd766_1 
+CB@6_mAd766_2 CB@6_mAd767_1 CB@6_mAd767_2 CB@6_mAd771_1 CB@6_mAd771_2 CB@6_mAd772_1 CB@6_mAd772_2 CB@6_mAd773_1 CB@6_mAd773_2 CB@6_mAd774_1 CB@6_mAd774_2 CB@6_mAd775_1 CB@6_mAd775_2 CB@6_mAd776_1 CB@6_mAd776_2 CB@6_mAd777_1 CB@6_mAd777_2 CB@6_X0 CB@6_X1 CB@6_X10 CB@6_X11 CB@6_X12 CB@6_X13 CB@6_X2 CB@6_X3 CB@6_X4 CB@6_X5 CB@6_X6 CB@6_X7 CB@6_X8 CB@6_X9 CB@6_Y1 CB@6_Y10 CB@6_Y11 CB@6_Y12 CB@6_Y2 CB@6_Y3 CB@6_Y4 CB@6_Y5 CB@6_Y6 CB@6_Y7 CB@6_Y8 CB@6_Y9 CB@6_Z1 CB@6_Z10 CB@6_Z11 CB@6_Z12 CB@6_Z2 CB@6_Z3 CB@6_Z4 
+CB@6_Z5 CB@6_Z6 CB@6_Z7 CB@6_Z8 CB@6_Z9 _5400TP094__CB
XCB@7 CB@7_K0 CB@7_K1 CB@7_K10 CB@7_K11 CB@7_K12 CB@7_K13 CB@7_K2 CB@7_K3 CB@7_K4 CB@7_K5 CB@7_K6 CB@7_K7 CB@7_K8 CB@7_K9 CB@7_mAd000_1 CB@7_mAd000_2 CB@7_mAd001_1 CB@7_mAd001_2 CB@7_mAd002_1 CB@7_mAd002_2 CB@7_mAd003_1 CB@7_mAd003_2 CB@7_mAd004_1 CB@7_mAd004_2 CB@7_mAd005_1 CB@7_mAd005_2 CB@7_mAd006_1 CB@7_mAd006_2 CB@7_mAd007_1 CB@7_mAd007_2 CB@7_mAd010_1 CB@7_mAd010_2 CB@7_mAd011_1 CB@7_mAd011_2 CB@7_mAd012_1 CB@7_mAd012_2 CB@7_mAd013_1 CB@7_mAd013_2 CB@7_mAd014_1 CB@7_mAd014_2 CB@7_mAd015_1 
+CB@7_mAd015_2 CB@7_mAd016_1 CB@7_mAd016_2 CB@7_mAd017_1 CB@7_mAd017_2 CB@7_mAd020_1 CB@7_mAd020_2 CB@7_mAd021_1 CB@7_mAd021_2 CB@7_mAd022_1 CB@7_mAd022_2 CB@7_mAd023_1 CB@7_mAd023_2 CB@7_mAd024_1 CB@7_mAd024_2 CB@7_mAd025_1 CB@7_mAd025_2 CB@7_mAd026_1 CB@7_mAd026_2 CB@7_mAd027_1 CB@7_mAd027_2 CB@7_mAd030_1 CB@7_mAd030_2 CB@7_mAd031_1 CB@7_mAd031_2 CB@7_mAd032_1 CB@7_mAd032_2 CB@7_mAd033_1 CB@7_mAd033_2 CB@7_mAd034_1 CB@7_mAd034_2 CB@7_mAd035_1 CB@7_mAd035_2 CB@7_mAd036_1 CB@7_mAd036_2 CB@7_mAd037_1 
+CB@7_mAd037_2 CB@7_mAd040_1 CB@7_mAd040_2 CB@7_mAd041_1 CB@7_mAd041_2 CB@7_mAd042_1 CB@7_mAd042_2 CB@7_mAd043_1 CB@7_mAd043_2 CB@7_mAd044_1 CB@7_mAd044_2 CB@7_mAd045_1 CB@7_mAd045_2 CB@7_mAd046_1 CB@7_mAd046_2 CB@7_mAd047_1 CB@7_mAd047_2 CB@7_mAd050_1 CB@7_mAd050_2 CB@7_mAd051_1 CB@7_mAd051_2 CB@7_mAd052_1 CB@7_mAd052_2 CB@7_mAd053_1 CB@7_mAd053_2 CB@7_mAd054_1 CB@7_mAd054_2 CB@7_mAd055_1 CB@7_mAd055_2 CB@7_mAd056_1 CB@7_mAd056_2 CB@7_mAd057_1 CB@7_mAd057_2 CB@7_mAd060_1 CB@7_mAd060_2 CB@7_mAd066_1 
+CB@7_mAd066_2 CB@7_mAd067_1 CB@7_mAd067_2 CB@7_mAd100_1 CB@7_mAd100_2 CB@7_mAd101_1 CB@7_mAd101_2 CB@7_mAd102_1 CB@7_mAd102_2 CB@7_mAd110_1 CB@7_mAd110_2 CB@7_mAd111_1 CB@7_mAd111_2 CB@7_mAd112_1 CB@7_mAd112_2 CB@7_mAd113_1 CB@7_mAd113_2 CB@7_mAd114_1 CB@7_mAd114_2 CB@7_mAd115_1 CB@7_mAd115_2 CB@7_mAd116_1 CB@7_mAd116_2 CB@7_mAd117_1 CB@7_mAd117_2 CB@7_mAd120_1 CB@7_mAd120_2 CB@7_mAd121_1 CB@7_mAd121_2 CB@7_mAd122_1 CB@7_mAd122_2 CB@7_mAd123_1 CB@7_mAd123_2 CB@7_mAd124_1 CB@7_mAd124_2 CB@7_mAd125_1 
+CB@7_mAd125_2 CB@7_mAd126_1 CB@7_mAd126_2 CB@7_mAd127_1 CB@7_mAd127_2 CB@7_mAd130_1 CB@7_mAd130_2 CB@7_mAd131_1 CB@7_mAd131_2 CB@7_mAd132_1 CB@7_mAd132_2 CB@7_mAd133_1 CB@7_mAd133_2 CB@7_mAd134_1 CB@7_mAd134_2 CB@7_mAd135_1 CB@7_mAd135_2 CB@7_mAd136_1 CB@7_mAd136_2 CB@7_mAd137_1 CB@7_mAd137_2 CB@7_mAd140_1 CB@7_mAd140_2 CB@7_mAd141_1 CB@7_mAd141_2 CB@7_mAd142_1 CB@7_mAd142_2 CB@7_mAd143_1 CB@7_mAd143_2 CB@7_mAd144_1 CB@7_mAd144_2 CB@7_mAd145_1 CB@7_mAd145_2 CB@7_mAd146_1 CB@7_mAd146_2 CB@7_mAd147_1 
+CB@7_mAd147_2 CB@7_mAd150_1 CB@7_mAd150_2 CB@7_mAd151_1 CB@7_mAd151_2 CB@7_mAd152_1 CB@7_mAd152_2 CB@7_mAd153_1 CB@7_mAd153_2 CB@7_mAd154_1 CB@7_mAd154_2 CB@7_mAd155_1 CB@7_mAd155_2 CB@7_mAd156_1 CB@7_mAd156_2 CB@7_mAd157_1 CB@7_mAd157_2 CB@7_mAd160_1 CB@7_mAd160_2 CB@7_mAd161_1 CB@7_mAd161_2 CB@7_mAd162_1 CB@7_mAd162_2 CB@7_mAd163_1 CB@7_mAd163_2 CB@7_mAd164_1 CB@7_mAd164_2 CB@7_mAd165_1 CB@7_mAd165_2 CB@7_mAd166_1 CB@7_mAd166_2 CB@7_mAd167_1 CB@7_mAd167_2 CB@7_mAd170_1 CB@7_mAd170_2 CB@7_mAd171_1 
+CB@7_mAd171_2 CB@7_mAd172_1 CB@7_mAd172_2 CB@7_mAd173_1 CB@7_mAd173_2 CB@7_mAd175_1 CB@7_mAd175_2 CB@7_mAd176_1 CB@7_mAd176_2 CB@7_mAd177_1 CB@7_mAd177_2 CB@7_mAd200_1 CB@7_mAd200_2 CB@7_mAd201_1 CB@7_mAd201_2 CB@7_mAd202_1 CB@7_mAd202_2 CB@7_mAd204_1 CB@7_mAd204_2 CB@7_mAd205_1 CB@7_mAd205_2 CB@7_mAd206_1 CB@7_mAd206_2 CB@7_mAd207_1 CB@7_mAd207_2 CB@7_mAd210_1 CB@7_mAd210_2 CB@7_mAd211_1 CB@7_mAd211_2 CB@7_mAd212_1 CB@7_mAd212_2 CB@7_mAd213_1 CB@7_mAd213_2 CB@7_mAd214_1 CB@7_mAd214_2 CB@7_mAd215_1 
+CB@7_mAd215_2 CB@7_mAd216_1 CB@7_mAd216_2 CB@7_mAd217_1 CB@7_mAd217_2 CB@7_mAd220_1 CB@7_mAd220_2 CB@7_mAd221_1 CB@7_mAd221_2 CB@7_mAd222_1 CB@7_mAd222_2 CB@7_mAd223_1 CB@7_mAd223_2 CB@7_mAd224_1 CB@7_mAd224_2 CB@7_mAd225_1 CB@7_mAd225_2 CB@7_mAd226_1 CB@7_mAd226_2 CB@7_mAd227_1 CB@7_mAd227_2 CB@7_mAd230_1 CB@7_mAd230_2 CB@7_mAd231_1 CB@7_mAd231_2 CB@7_mAd232_1 CB@7_mAd232_2 CB@7_mAd233_1 CB@7_mAd233_2 CB@7_mAd234_1 CB@7_mAd234_2 CB@7_mAd235_1 CB@7_mAd235_2 CB@7_mAd236_1 CB@7_mAd236_2 CB@7_mAd237_1 
+CB@7_mAd237_2 CB@7_mAd240_1 CB@7_mAd240_2 CB@7_mAd241_1 CB@7_mAd241_2 CB@7_mAd242_1 CB@7_mAd242_2 CB@7_mAd243_1 CB@7_mAd243_2 CB@7_mAd244_1 CB@7_mAd244_2 CB@7_mAd245_1 CB@7_mAd245_2 CB@7_mAd246_1 CB@7_mAd246_2 CB@7_mAd247_1 CB@7_mAd247_2 CB@7_mAd250_1 CB@7_mAd250_2 CB@7_mAd251_1 CB@7_mAd251_2 CB@7_mAd252_1 CB@7_mAd252_2 CB@7_mAd253_1 CB@7_mAd253_2 CB@7_mAd254_1 CB@7_mAd254_2 CB@7_mAd255_1 CB@7_mAd255_2 CB@7_mAd256_1 CB@7_mAd256_2 CB@7_mAd257_1 CB@7_mAd257_2 CB@7_mAd260_1 CB@7_mAd260_2 CB@7_mAd261_1 
+CB@7_mAd261_2 CB@7_mAd262_1 CB@7_mAd262_2 CB@7_mAd263_1 CB@7_mAd263_2 CB@7_mAd264_1 CB@7_mAd264_2 CB@7_mAd265_1 CB@7_mAd265_2 CB@7_mAd266_1 CB@7_mAd266_2 CB@7_mAd267_1 CB@7_mAd267_2 CB@7_mAd275_1 CB@7_mAd275_2 CB@7_mAd276_1 CB@7_mAd276_2 CB@7_mAd277_1 CB@7_mAd277_2 CB@7_mAd300_1 CB@7_mAd300_2 CB@7_mAd310_1 CB@7_mAd310_2 CB@7_mAd311_1 CB@7_mAd311_2 CB@7_mAd317_1 CB@7_mAd317_2 CB@7_mAd320_1 CB@7_mAd320_2 CB@7_mAd321_1 CB@7_mAd321_2 CB@7_mAd322_1 CB@7_mAd322_2 CB@7_mAd323_1 CB@7_mAd323_2 CB@7_mAd324_1 
+CB@7_mAd324_2 CB@7_mAd325_1 CB@7_mAd325_2 CB@7_mAd326_1 CB@7_mAd326_2 CB@7_mAd327_1 CB@7_mAd327_2 CB@7_mAd330_1 CB@7_mAd330_2 CB@7_mAd331_1 CB@7_mAd331_2 CB@7_mAd332_1 CB@7_mAd332_2 CB@7_mAd333_1 CB@7_mAd333_2 CB@7_mAd334_1 CB@7_mAd334_2 CB@7_mAd335_1 CB@7_mAd335_2 CB@7_mAd336_1 CB@7_mAd336_2 CB@7_mAd337_1 CB@7_mAd337_2 CB@7_mAd340_1 CB@7_mAd340_2 CB@7_mAd341_1 CB@7_mAd341_2 CB@7_mAd342_1 CB@7_mAd342_2 CB@7_mAd343_1 CB@7_mAd343_2 CB@7_mAd344_1 CB@7_mAd344_2 CB@7_mAd345_1 CB@7_mAd345_2 CB@7_mAd346_1 
+CB@7_mAd346_2 CB@7_mAd347_1 CB@7_mAd347_2 CB@7_mAd350_1 CB@7_mAd350_2 CB@7_mAd351_1 CB@7_mAd351_2 CB@7_mAd352_1 CB@7_mAd352_2 CB@7_mAd353_1 CB@7_mAd353_2 CB@7_mAd354_1 CB@7_mAd354_2 CB@7_mAd355_1 CB@7_mAd355_2 CB@7_mAd356_1 CB@7_mAd356_2 CB@7_mAd357_1 CB@7_mAd357_2 CB@7_mAd360_1 CB@7_mAd360_2 CB@7_mAd361_1 CB@7_mAd361_2 CB@7_mAd362_1 CB@7_mAd362_2 CB@7_mAd363_1 CB@7_mAd363_2 CB@7_mAd364_1 CB@7_mAd364_2 CB@7_mAd365_1 CB@7_mAd365_2 CB@7_mAd366_1 CB@7_mAd366_2 CB@7_mAd367_1 CB@7_mAd367_2 CB@7_mAd371_1 
+CB@7_mAd371_2 CB@7_mAd372_1 CB@7_mAd372_2 CB@7_mAd373_1 CB@7_mAd373_2 CB@7_mAd374_1 CB@7_mAd374_2 CB@7_mAd375_1 CB@7_mAd375_2 CB@7_mAd376_1 CB@7_mAd376_2 CB@7_mAd377_1 CB@7_mAd377_2 CB@7_mAd400_1 CB@7_mAd400_2 CB@7_mAd401_1 CB@7_mAd401_2 CB@7_mAd402_1 CB@7_mAd402_2 CB@7_mAd403_1 CB@7_mAd403_2 CB@7_mAd404_1 CB@7_mAd404_2 CB@7_mAd405_1 CB@7_mAd405_2 CB@7_mAd406_1 CB@7_mAd406_2 CB@7_mAd407_1 CB@7_mAd407_2 CB@7_mAd410_1 CB@7_mAd410_2 CB@7_mAd411_1 CB@7_mAd411_2 CB@7_mAd412_1 CB@7_mAd412_2 CB@7_mAd413_1 
+CB@7_mAd413_2 CB@7_mAd414_1 CB@7_mAd414_2 CB@7_mAd415_1 CB@7_mAd415_2 CB@7_mAd416_1 CB@7_mAd416_2 CB@7_mAd417_1 CB@7_mAd417_2 CB@7_mAd420_1 CB@7_mAd420_2 CB@7_mAd421_1 CB@7_mAd421_2 CB@7_mAd422_1 CB@7_mAd422_2 CB@7_mAd423_1 CB@7_mAd423_2 CB@7_mAd424_1 CB@7_mAd424_2 CB@7_mAd425_1 CB@7_mAd425_2 CB@7_mAd426_1 CB@7_mAd426_2 CB@7_mAd427_1 CB@7_mAd427_2 CB@7_mAd430_1 CB@7_mAd430_2 CB@7_mAd431_1 CB@7_mAd431_2 CB@7_mAd432_1 CB@7_mAd432_2 CB@7_mAd433_1 CB@7_mAd433_2 CB@7_mAd434_1 CB@7_mAd434_2 CB@7_mAd435_1 
+CB@7_mAd435_2 CB@7_mAd436_1 CB@7_mAd436_2 CB@7_mAd437_1 CB@7_mAd437_2 CB@7_mAd440_1 CB@7_mAd440_2 CB@7_mAd441_1 CB@7_mAd441_2 CB@7_mAd442_1 CB@7_mAd442_2 CB@7_mAd443_1 CB@7_mAd443_2 CB@7_mAd444_1 CB@7_mAd444_2 CB@7_mAd445_1 CB@7_mAd445_2 CB@7_mAd446_1 CB@7_mAd446_2 CB@7_mAd447_1 CB@7_mAd447_2 CB@7_mAd450_1 CB@7_mAd450_2 CB@7_mAd451_1 CB@7_mAd451_2 CB@7_mAd452_1 CB@7_mAd452_2 CB@7_mAd453_1 CB@7_mAd453_2 CB@7_mAd454_1 CB@7_mAd454_2 CB@7_mAd455_1 CB@7_mAd455_2 CB@7_mAd456_1 CB@7_mAd456_2 CB@7_mAd457_1 
+CB@7_mAd457_2 CB@7_mAd460_1 CB@7_mAd460_2 CB@7_mAd466_1 CB@7_mAd466_2 CB@7_mAd467_1 CB@7_mAd467_2 CB@7_mAd500_1 CB@7_mAd500_2 CB@7_mAd501_1 CB@7_mAd501_2 CB@7_mAd502_1 CB@7_mAd502_2 CB@7_mAd508_1 CB@7_mAd508_2 CB@7_mAd509_1 CB@7_mAd509_2 CB@7_mAd512_1 CB@7_mAd512_2 CB@7_mAd513_1 CB@7_mAd513_2 CB@7_mAd514_1 CB@7_mAd514_2 CB@7_mAd515_1 CB@7_mAd515_2 CB@7_mAd516_1 CB@7_mAd516_2 CB@7_mAd517_1 CB@7_mAd517_2 CB@7_mAd520_1 CB@7_mAd520_2 CB@7_mAd521_1 CB@7_mAd521_2 CB@7_mAd522_1 CB@7_mAd522_2 CB@7_mAd523_1 
+CB@7_mAd523_2 CB@7_mAd524_1 CB@7_mAd524_2 CB@7_mAd525_1 CB@7_mAd525_2 CB@7_mAd526_1 CB@7_mAd526_2 CB@7_mAd527_1 CB@7_mAd527_2 CB@7_mAd530_1 CB@7_mAd530_2 CB@7_mAd531_1 CB@7_mAd531_2 CB@7_mAd532_1 CB@7_mAd532_2 CB@7_mAd533_1 CB@7_mAd533_2 CB@7_mAd534_1 CB@7_mAd534_2 CB@7_mAd535_1 CB@7_mAd535_2 CB@7_mAd536_1 CB@7_mAd536_2 CB@7_mAd537_1 CB@7_mAd537_2 CB@7_mAd540_1 CB@7_mAd540_2 CB@7_mAd541_1 CB@7_mAd541_2 CB@7_mAd542_1 CB@7_mAd542_2 CB@7_mAd543_1 CB@7_mAd543_2 CB@7_mAd544_1 CB@7_mAd544_2 CB@7_mAd545_1 
+CB@7_mAd545_2 CB@7_mAd546_1 CB@7_mAd546_2 CB@7_mAd547_1 CB@7_mAd547_2 CB@7_mAd550_1 CB@7_mAd550_2 CB@7_mAd551_1 CB@7_mAd551_2 CB@7_mAd552_1 CB@7_mAd552_2 CB@7_mAd553_1 CB@7_mAd553_2 CB@7_mAd554_1 CB@7_mAd554_2 CB@7_mAd555_1 CB@7_mAd555_2 CB@7_mAd556_1 CB@7_mAd556_2 CB@7_mAd557_1 CB@7_mAd557_2 CB@7_mAd560_1 CB@7_mAd560_2 CB@7_mAd561_1 CB@7_mAd561_2 CB@7_mAd562_1 CB@7_mAd562_2 CB@7_mAd563_1 CB@7_mAd563_2 CB@7_mAd564_1 CB@7_mAd564_2 CB@7_mAd565_1 CB@7_mAd565_2 CB@7_mAd566_1 CB@7_mAd566_2 CB@7_mAd567_1 
+CB@7_mAd567_2 CB@7_mAd570_1 CB@7_mAd570_2 CB@7_mAd571_1 CB@7_mAd571_2 CB@7_mAd572_1 CB@7_mAd572_2 CB@7_mAd573_1 CB@7_mAd573_2 CB@7_mAd575_1 CB@7_mAd575_2 CB@7_mAd576_1 CB@7_mAd576_2 CB@7_mAd577_1 CB@7_mAd577_2 CB@7_mAd600_1 CB@7_mAd600_2 CB@7_mAd601_1 CB@7_mAd601_2 CB@7_mAd602_1 CB@7_mAd602_2 CB@7_mAd604_1 CB@7_mAd604_2 CB@7_mAd605_1 CB@7_mAd605_2 CB@7_mAd606_1 CB@7_mAd606_2 CB@7_mAd607_1 CB@7_mAd607_2 CB@7_mAd610_1 CB@7_mAd610_2 CB@7_mAd611_1 CB@7_mAd611_2 CB@7_mAd612_1 CB@7_mAd612_2 CB@7_mAd613_1 
+CB@7_mAd613_2 CB@7_mAd614_1 CB@7_mAd614_2 CB@7_mAd615_1 CB@7_mAd615_2 CB@7_mAd616_1 CB@7_mAd616_2 CB@7_mAd617_1 CB@7_mAd617_2 CB@7_mAd620_1 CB@7_mAd620_2 CB@7_mAd621_1 CB@7_mAd621_2 CB@7_mAd622_1 CB@7_mAd622_2 CB@7_mAd623_1 CB@7_mAd623_2 CB@7_mAd624_1 CB@7_mAd624_2 CB@7_mAd625_1 CB@7_mAd625_2 CB@7_mAd626_1 CB@7_mAd626_2 CB@7_mAd627_1 CB@7_mAd627_2 CB@7_mAd630_1 CB@7_mAd630_2 CB@7_mAd631_1 CB@7_mAd631_2 CB@7_mAd632_1 CB@7_mAd632_2 CB@7_mAd633_1 CB@7_mAd633_2 CB@7_mAd634_1 CB@7_mAd634_2 CB@7_mAd635_1 
+CB@7_mAd635_2 CB@7_mAd636_1 CB@7_mAd636_2 CB@7_mAd637_1 CB@7_mAd637_2 CB@7_mAd640_1 CB@7_mAd640_2 CB@7_mAd641_1 CB@7_mAd641_2 CB@7_mAd642_1 CB@7_mAd642_2 CB@7_mAd643_1 CB@7_mAd643_2 CB@7_mAd644_1 CB@7_mAd644_2 CB@7_mAd645_1 CB@7_mAd645_2 CB@7_mAd646_1 CB@7_mAd646_2 CB@7_mAd647_1 CB@7_mAd647_2 CB@7_mAd650_1 CB@7_mAd650_2 CB@7_mAd651_1 CB@7_mAd651_2 CB@7_mAd652_1 CB@7_mAd652_2 CB@7_mAd653_1 CB@7_mAd653_2 CB@7_mAd654_1 CB@7_mAd654_2 CB@7_mAd655_1 CB@7_mAd655_2 CB@7_mAd656_1 CB@7_mAd656_2 CB@7_mAd657_1 
+CB@7_mAd657_2 CB@7_mAd660_1 CB@7_mAd660_2 CB@7_mAd661_1 CB@7_mAd661_2 CB@7_mAd662_1 CB@7_mAd662_2 CB@7_mAd663_1 CB@7_mAd663_2 CB@7_mAd664_1 CB@7_mAd664_2 CB@7_mAd665_1 CB@7_mAd665_2 CB@7_mAd666_1 CB@7_mAd666_2 CB@7_mAd667_1 CB@7_mAd667_2 CB@7_mAd675_1 CB@7_mAd675_2 CB@7_mAd676_1 CB@7_mAd676_2 CB@7_mAd677_1 CB@7_mAd677_2 CB@7_mAd700_1 CB@7_mAd700_2 CB@7_mAd710_1 CB@7_mAd710_2 CB@7_mAd711_1 CB@7_mAd711_2 CB@7_mAd717_1 CB@7_mAd717_2 CB@7_mAd720_1 CB@7_mAd720_2 CB@7_mAd721_1 CB@7_mAd721_2 CB@7_mAd722_1 
+CB@7_mAd722_2 CB@7_mAd723_1 CB@7_mAd723_2 CB@7_mAd724_1 CB@7_mAd724_2 CB@7_mAd725_1 CB@7_mAd725_2 CB@7_mAd726_1 CB@7_mAd726_2 CB@7_mAd727_1 CB@7_mAd727_2 CB@7_mAd730_1 CB@7_mAd730_2 CB@7_mAd731_1 CB@7_mAd731_2 CB@7_mAd732_1 CB@7_mAd732_2 CB@7_mAd733_1 CB@7_mAd733_2 CB@7_mAd734_1 CB@7_mAd734_2 CB@7_mAd735_1 CB@7_mAd735_2 CB@7_mAd736_1 CB@7_mAd736_2 CB@7_mAd737_1 CB@7_mAd737_2 CB@7_mAd740_1 CB@7_mAd740_2 CB@7_mAd741_1 CB@7_mAd741_2 CB@7_mAd742_1 CB@7_mAd742_2 CB@7_mAd743_1 CB@7_mAd743_2 CB@7_mAd744_1 
+CB@7_mAd744_2 CB@7_mAd745_1 CB@7_mAd745_2 CB@7_mAd746_1 CB@7_mAd746_2 CB@7_mAd747_1 CB@7_mAd747_2 CB@7_mAd750_1 CB@7_mAd750_2 CB@7_mAd751_1 CB@7_mAd751_2 CB@7_mAd752_1 CB@7_mAd752_2 CB@7_mAd753_1 CB@7_mAd753_2 CB@7_mAd754_1 CB@7_mAd754_2 CB@7_mAd755_1 CB@7_mAd755_2 CB@7_mAd756_1 CB@7_mAd756_2 CB@7_mAd757_1 CB@7_mAd757_2 CB@7_mAd760_1 CB@7_mAd760_2 CB@7_mAd761_1 CB@7_mAd761_2 CB@7_mAd762_1 CB@7_mAd762_2 CB@7_mAd763_1 CB@7_mAd763_2 CB@7_mAd764_1 CB@7_mAd764_2 CB@7_mAd765_1 CB@7_mAd765_2 CB@7_mAd766_1 
+CB@7_mAd766_2 CB@7_mAd767_1 CB@7_mAd767_2 CB@7_mAd771_1 CB@7_mAd771_2 CB@7_mAd772_1 CB@7_mAd772_2 CB@7_mAd773_1 CB@7_mAd773_2 CB@7_mAd774_1 CB@7_mAd774_2 CB@7_mAd775_1 CB@7_mAd775_2 CB@7_mAd776_1 CB@7_mAd776_2 CB@7_mAd777_1 CB@7_mAd777_2 CB@7_X0 CB@7_X1 CB@7_X10 CB@7_X11 CB@7_X12 CB@7_X13 CB@7_X2 CB@7_X3 CB@7_X4 CB@7_X5 CB@7_X6 CB@7_X7 CB@7_X8 CB@7_X9 CB@7_Y1 CB@7_Y10 CB@7_Y11 CB@7_Y12 CB@7_Y2 CB@7_Y3 CB@7_Y4 CB@7_Y5 CB@7_Y6 CB@7_Y7 CB@7_Y8 CB@7_Y9 CB@7_Z1 CB@7_Z10 CB@7_Z11 CB@7_Z12 CB@7_Z2 CB@7_Z3 CB@7_Z4 
+CB@7_Z5 CB@7_Z6 CB@7_Z7 CB@7_Z8 CB@7_Z9 _5400TP094__CB
XCB@8 CB@8_K0 CB@8_K1 CB@8_K10 CB@8_K11 CB@8_K12 CB@8_K13 CB@8_K2 CB@8_K3 CB@8_K4 CB@8_K5 CB@8_K6 CB@8_K7 CB@8_K8 CB@8_K9 CB@8_mAd000_1 CB@8_mAd000_2 CB@8_mAd001_1 CB@8_mAd001_2 CB@8_mAd002_1 CB@8_mAd002_2 CB@8_mAd003_1 CB@8_mAd003_2 CB@8_mAd004_1 CB@8_mAd004_2 CB@8_mAd005_1 CB@8_mAd005_2 CB@8_mAd006_1 CB@8_mAd006_2 CB@8_mAd007_1 CB@8_mAd007_2 CB@8_mAd010_1 CB@8_mAd010_2 CB@8_mAd011_1 CB@8_mAd011_2 CB@8_mAd012_1 CB@8_mAd012_2 CB@8_mAd013_1 CB@8_mAd013_2 CB@8_mAd014_1 CB@8_mAd014_2 CB@8_mAd015_1 
+CB@8_mAd015_2 CB@8_mAd016_1 CB@8_mAd016_2 CB@8_mAd017_1 CB@8_mAd017_2 CB@8_mAd020_1 CB@8_mAd020_2 CB@8_mAd021_1 CB@8_mAd021_2 CB@8_mAd022_1 CB@8_mAd022_2 CB@8_mAd023_1 CB@8_mAd023_2 CB@8_mAd024_1 CB@8_mAd024_2 CB@8_mAd025_1 CB@8_mAd025_2 CB@8_mAd026_1 CB@8_mAd026_2 CB@8_mAd027_1 CB@8_mAd027_2 CB@8_mAd030_1 CB@8_mAd030_2 CB@8_mAd031_1 CB@8_mAd031_2 CB@8_mAd032_1 CB@8_mAd032_2 CB@8_mAd033_1 CB@8_mAd033_2 CB@8_mAd034_1 CB@8_mAd034_2 CB@8_mAd035_1 CB@8_mAd035_2 CB@8_mAd036_1 CB@8_mAd036_2 CB@8_mAd037_1 
+CB@8_mAd037_2 CB@8_mAd040_1 CB@8_mAd040_2 CB@8_mAd041_1 CB@8_mAd041_2 CB@8_mAd042_1 CB@8_mAd042_2 CB@8_mAd043_1 CB@8_mAd043_2 CB@8_mAd044_1 CB@8_mAd044_2 CB@8_mAd045_1 CB@8_mAd045_2 CB@8_mAd046_1 CB@8_mAd046_2 CB@8_mAd047_1 CB@8_mAd047_2 CB@8_mAd050_1 CB@8_mAd050_2 CB@8_mAd051_1 CB@8_mAd051_2 CB@8_mAd052_1 CB@8_mAd052_2 CB@8_mAd053_1 CB@8_mAd053_2 CB@8_mAd054_1 CB@8_mAd054_2 CB@8_mAd055_1 CB@8_mAd055_2 CB@8_mAd056_1 CB@8_mAd056_2 CB@8_mAd057_1 CB@8_mAd057_2 CB@8_mAd060_1 CB@8_mAd060_2 CB@8_mAd066_1 
+CB@8_mAd066_2 CB@8_mAd067_1 CB@8_mAd067_2 CB@8_mAd100_1 CB@8_mAd100_2 CB@8_mAd101_1 CB@8_mAd101_2 CB@8_mAd102_1 CB@8_mAd102_2 CB@8_mAd110_1 CB@8_mAd110_2 CB@8_mAd111_1 CB@8_mAd111_2 CB@8_mAd112_1 CB@8_mAd112_2 CB@8_mAd113_1 CB@8_mAd113_2 CB@8_mAd114_1 CB@8_mAd114_2 CB@8_mAd115_1 CB@8_mAd115_2 CB@8_mAd116_1 CB@8_mAd116_2 CB@8_mAd117_1 CB@8_mAd117_2 CB@8_mAd120_1 CB@8_mAd120_2 CB@8_mAd121_1 CB@8_mAd121_2 CB@8_mAd122_1 CB@8_mAd122_2 CB@8_mAd123_1 CB@8_mAd123_2 CB@8_mAd124_1 CB@8_mAd124_2 CB@8_mAd125_1 
+CB@8_mAd125_2 CB@8_mAd126_1 CB@8_mAd126_2 CB@8_mAd127_1 CB@8_mAd127_2 CB@8_mAd130_1 CB@8_mAd130_2 CB@8_mAd131_1 CB@8_mAd131_2 CB@8_mAd132_1 CB@8_mAd132_2 CB@8_mAd133_1 CB@8_mAd133_2 CB@8_mAd134_1 CB@8_mAd134_2 CB@8_mAd135_1 CB@8_mAd135_2 CB@8_mAd136_1 CB@8_mAd136_2 CB@8_mAd137_1 CB@8_mAd137_2 CB@8_mAd140_1 CB@8_mAd140_2 CB@8_mAd141_1 CB@8_mAd141_2 CB@8_mAd142_1 CB@8_mAd142_2 CB@8_mAd143_1 CB@8_mAd143_2 CB@8_mAd144_1 CB@8_mAd144_2 CB@8_mAd145_1 CB@8_mAd145_2 CB@8_mAd146_1 CB@8_mAd146_2 CB@8_mAd147_1 
+CB@8_mAd147_2 CB@8_mAd150_1 CB@8_mAd150_2 CB@8_mAd151_1 CB@8_mAd151_2 CB@8_mAd152_1 CB@8_mAd152_2 CB@8_mAd153_1 CB@8_mAd153_2 CB@8_mAd154_1 CB@8_mAd154_2 CB@8_mAd155_1 CB@8_mAd155_2 CB@8_mAd156_1 CB@8_mAd156_2 CB@8_mAd157_1 CB@8_mAd157_2 CB@8_mAd160_1 CB@8_mAd160_2 CB@8_mAd161_1 CB@8_mAd161_2 CB@8_mAd162_1 CB@8_mAd162_2 CB@8_mAd163_1 CB@8_mAd163_2 CB@8_mAd164_1 CB@8_mAd164_2 CB@8_mAd165_1 CB@8_mAd165_2 CB@8_mAd166_1 CB@8_mAd166_2 CB@8_mAd167_1 CB@8_mAd167_2 CB@8_mAd170_1 CB@8_mAd170_2 CB@8_mAd171_1 
+CB@8_mAd171_2 CB@8_mAd172_1 CB@8_mAd172_2 CB@8_mAd173_1 CB@8_mAd173_2 CB@8_mAd175_1 CB@8_mAd175_2 CB@8_mAd176_1 CB@8_mAd176_2 CB@8_mAd177_1 CB@8_mAd177_2 CB@8_mAd200_1 CB@8_mAd200_2 CB@8_mAd201_1 CB@8_mAd201_2 CB@8_mAd202_1 CB@8_mAd202_2 CB@8_mAd204_1 CB@8_mAd204_2 CB@8_mAd205_1 CB@8_mAd205_2 CB@8_mAd206_1 CB@8_mAd206_2 CB@8_mAd207_1 CB@8_mAd207_2 CB@8_mAd210_1 CB@8_mAd210_2 CB@8_mAd211_1 CB@8_mAd211_2 CB@8_mAd212_1 CB@8_mAd212_2 CB@8_mAd213_1 CB@8_mAd213_2 CB@8_mAd214_1 CB@8_mAd214_2 CB@8_mAd215_1 
+CB@8_mAd215_2 CB@8_mAd216_1 CB@8_mAd216_2 CB@8_mAd217_1 CB@8_mAd217_2 CB@8_mAd220_1 CB@8_mAd220_2 CB@8_mAd221_1 CB@8_mAd221_2 CB@8_mAd222_1 CB@8_mAd222_2 CB@8_mAd223_1 CB@8_mAd223_2 CB@8_mAd224_1 CB@8_mAd224_2 CB@8_mAd225_1 CB@8_mAd225_2 CB@8_mAd226_1 CB@8_mAd226_2 CB@8_mAd227_1 CB@8_mAd227_2 CB@8_mAd230_1 CB@8_mAd230_2 CB@8_mAd231_1 CB@8_mAd231_2 CB@8_mAd232_1 CB@8_mAd232_2 CB@8_mAd233_1 CB@8_mAd233_2 CB@8_mAd234_1 CB@8_mAd234_2 CB@8_mAd235_1 CB@8_mAd235_2 CB@8_mAd236_1 CB@8_mAd236_2 CB@8_mAd237_1 
+CB@8_mAd237_2 CB@8_mAd240_1 CB@8_mAd240_2 CB@8_mAd241_1 CB@8_mAd241_2 CB@8_mAd242_1 CB@8_mAd242_2 CB@8_mAd243_1 CB@8_mAd243_2 CB@8_mAd244_1 CB@8_mAd244_2 CB@8_mAd245_1 CB@8_mAd245_2 CB@8_mAd246_1 CB@8_mAd246_2 CB@8_mAd247_1 CB@8_mAd247_2 CB@8_mAd250_1 CB@8_mAd250_2 CB@8_mAd251_1 CB@8_mAd251_2 CB@8_mAd252_1 CB@8_mAd252_2 CB@8_mAd253_1 CB@8_mAd253_2 CB@8_mAd254_1 CB@8_mAd254_2 CB@8_mAd255_1 CB@8_mAd255_2 CB@8_mAd256_1 CB@8_mAd256_2 CB@8_mAd257_1 CB@8_mAd257_2 CB@8_mAd260_1 CB@8_mAd260_2 CB@8_mAd261_1 
+CB@8_mAd261_2 CB@8_mAd262_1 CB@8_mAd262_2 CB@8_mAd263_1 CB@8_mAd263_2 CB@8_mAd264_1 CB@8_mAd264_2 CB@8_mAd265_1 CB@8_mAd265_2 CB@8_mAd266_1 CB@8_mAd266_2 CB@8_mAd267_1 CB@8_mAd267_2 CB@8_mAd275_1 CB@8_mAd275_2 CB@8_mAd276_1 CB@8_mAd276_2 CB@8_mAd277_1 CB@8_mAd277_2 CB@8_mAd300_1 CB@8_mAd300_2 CB@8_mAd310_1 CB@8_mAd310_2 CB@8_mAd311_1 CB@8_mAd311_2 CB@8_mAd317_1 CB@8_mAd317_2 CB@8_mAd320_1 CB@8_mAd320_2 CB@8_mAd321_1 CB@8_mAd321_2 CB@8_mAd322_1 CB@8_mAd322_2 CB@8_mAd323_1 CB@8_mAd323_2 CB@8_mAd324_1 
+CB@8_mAd324_2 CB@8_mAd325_1 CB@8_mAd325_2 CB@8_mAd326_1 CB@8_mAd326_2 CB@8_mAd327_1 CB@8_mAd327_2 CB@8_mAd330_1 CB@8_mAd330_2 CB@8_mAd331_1 CB@8_mAd331_2 CB@8_mAd332_1 CB@8_mAd332_2 CB@8_mAd333_1 CB@8_mAd333_2 CB@8_mAd334_1 CB@8_mAd334_2 CB@8_mAd335_1 CB@8_mAd335_2 CB@8_mAd336_1 CB@8_mAd336_2 CB@8_mAd337_1 CB@8_mAd337_2 CB@8_mAd340_1 CB@8_mAd340_2 CB@8_mAd341_1 CB@8_mAd341_2 CB@8_mAd342_1 CB@8_mAd342_2 CB@8_mAd343_1 CB@8_mAd343_2 CB@8_mAd344_1 CB@8_mAd344_2 CB@8_mAd345_1 CB@8_mAd345_2 CB@8_mAd346_1 
+CB@8_mAd346_2 CB@8_mAd347_1 CB@8_mAd347_2 CB@8_mAd350_1 CB@8_mAd350_2 CB@8_mAd351_1 CB@8_mAd351_2 CB@8_mAd352_1 CB@8_mAd352_2 CB@8_mAd353_1 CB@8_mAd353_2 CB@8_mAd354_1 CB@8_mAd354_2 CB@8_mAd355_1 CB@8_mAd355_2 CB@8_mAd356_1 CB@8_mAd356_2 CB@8_mAd357_1 CB@8_mAd357_2 CB@8_mAd360_1 CB@8_mAd360_2 CB@8_mAd361_1 CB@8_mAd361_2 CB@8_mAd362_1 CB@8_mAd362_2 CB@8_mAd363_1 CB@8_mAd363_2 CB@8_mAd364_1 CB@8_mAd364_2 CB@8_mAd365_1 CB@8_mAd365_2 CB@8_mAd366_1 CB@8_mAd366_2 CB@8_mAd367_1 CB@8_mAd367_2 CB@8_mAd371_1 
+CB@8_mAd371_2 CB@8_mAd372_1 CB@8_mAd372_2 CB@8_mAd373_1 CB@8_mAd373_2 CB@8_mAd374_1 CB@8_mAd374_2 CB@8_mAd375_1 CB@8_mAd375_2 CB@8_mAd376_1 CB@8_mAd376_2 CB@8_mAd377_1 CB@8_mAd377_2 CB@8_mAd400_1 CB@8_mAd400_2 CB@8_mAd401_1 CB@8_mAd401_2 CB@8_mAd402_1 CB@8_mAd402_2 CB@8_mAd403_1 CB@8_mAd403_2 CB@8_mAd404_1 CB@8_mAd404_2 CB@8_mAd405_1 CB@8_mAd405_2 CB@8_mAd406_1 CB@8_mAd406_2 CB@8_mAd407_1 CB@8_mAd407_2 CB@8_mAd410_1 CB@8_mAd410_2 CB@8_mAd411_1 CB@8_mAd411_2 CB@8_mAd412_1 CB@8_mAd412_2 CB@8_mAd413_1 
+CB@8_mAd413_2 CB@8_mAd414_1 CB@8_mAd414_2 CB@8_mAd415_1 CB@8_mAd415_2 CB@8_mAd416_1 CB@8_mAd416_2 CB@8_mAd417_1 CB@8_mAd417_2 CB@8_mAd420_1 CB@8_mAd420_2 CB@8_mAd421_1 CB@8_mAd421_2 CB@8_mAd422_1 CB@8_mAd422_2 CB@8_mAd423_1 CB@8_mAd423_2 CB@8_mAd424_1 CB@8_mAd424_2 CB@8_mAd425_1 CB@8_mAd425_2 CB@8_mAd426_1 CB@8_mAd426_2 CB@8_mAd427_1 CB@8_mAd427_2 CB@8_mAd430_1 CB@8_mAd430_2 CB@8_mAd431_1 CB@8_mAd431_2 CB@8_mAd432_1 CB@8_mAd432_2 CB@8_mAd433_1 CB@8_mAd433_2 CB@8_mAd434_1 CB@8_mAd434_2 CB@8_mAd435_1 
+CB@8_mAd435_2 CB@8_mAd436_1 CB@8_mAd436_2 CB@8_mAd437_1 CB@8_mAd437_2 CB@8_mAd440_1 CB@8_mAd440_2 CB@8_mAd441_1 CB@8_mAd441_2 CB@8_mAd442_1 CB@8_mAd442_2 CB@8_mAd443_1 CB@8_mAd443_2 CB@8_mAd444_1 CB@8_mAd444_2 CB@8_mAd445_1 CB@8_mAd445_2 CB@8_mAd446_1 CB@8_mAd446_2 CB@8_mAd447_1 CB@8_mAd447_2 CB@8_mAd450_1 CB@8_mAd450_2 CB@8_mAd451_1 CB@8_mAd451_2 CB@8_mAd452_1 CB@8_mAd452_2 CB@8_mAd453_1 CB@8_mAd453_2 CB@8_mAd454_1 CB@8_mAd454_2 CB@8_mAd455_1 CB@8_mAd455_2 CB@8_mAd456_1 CB@8_mAd456_2 CB@8_mAd457_1 
+CB@8_mAd457_2 CB@8_mAd460_1 CB@8_mAd460_2 CB@8_mAd466_1 CB@8_mAd466_2 CB@8_mAd467_1 CB@8_mAd467_2 CB@8_mAd500_1 CB@8_mAd500_2 CB@8_mAd501_1 CB@8_mAd501_2 CB@8_mAd502_1 CB@8_mAd502_2 CB@8_mAd508_1 CB@8_mAd508_2 CB@8_mAd509_1 CB@8_mAd509_2 CB@8_mAd512_1 CB@8_mAd512_2 CB@8_mAd513_1 CB@8_mAd513_2 CB@8_mAd514_1 CB@8_mAd514_2 CB@8_mAd515_1 CB@8_mAd515_2 CB@8_mAd516_1 CB@8_mAd516_2 CB@8_mAd517_1 CB@8_mAd517_2 CB@8_mAd520_1 CB@8_mAd520_2 CB@8_mAd521_1 CB@8_mAd521_2 CB@8_mAd522_1 CB@8_mAd522_2 CB@8_mAd523_1 
+CB@8_mAd523_2 CB@8_mAd524_1 CB@8_mAd524_2 CB@8_mAd525_1 CB@8_mAd525_2 CB@8_mAd526_1 CB@8_mAd526_2 CB@8_mAd527_1 CB@8_mAd527_2 CB@8_mAd530_1 CB@8_mAd530_2 CB@8_mAd531_1 CB@8_mAd531_2 CB@8_mAd532_1 CB@8_mAd532_2 CB@8_mAd533_1 CB@8_mAd533_2 CB@8_mAd534_1 CB@8_mAd534_2 CB@8_mAd535_1 CB@8_mAd535_2 CB@8_mAd536_1 CB@8_mAd536_2 CB@8_mAd537_1 CB@8_mAd537_2 CB@8_mAd540_1 CB@8_mAd540_2 CB@8_mAd541_1 CB@8_mAd541_2 CB@8_mAd542_1 CB@8_mAd542_2 CB@8_mAd543_1 CB@8_mAd543_2 CB@8_mAd544_1 CB@8_mAd544_2 CB@8_mAd545_1 
+CB@8_mAd545_2 CB@8_mAd546_1 CB@8_mAd546_2 CB@8_mAd547_1 CB@8_mAd547_2 CB@8_mAd550_1 CB@8_mAd550_2 CB@8_mAd551_1 CB@8_mAd551_2 CB@8_mAd552_1 CB@8_mAd552_2 CB@8_mAd553_1 CB@8_mAd553_2 CB@8_mAd554_1 CB@8_mAd554_2 CB@8_mAd555_1 CB@8_mAd555_2 CB@8_mAd556_1 CB@8_mAd556_2 CB@8_mAd557_1 CB@8_mAd557_2 CB@8_mAd560_1 CB@8_mAd560_2 CB@8_mAd561_1 CB@8_mAd561_2 CB@8_mAd562_1 CB@8_mAd562_2 CB@8_mAd563_1 CB@8_mAd563_2 CB@8_mAd564_1 CB@8_mAd564_2 CB@8_mAd565_1 CB@8_mAd565_2 CB@8_mAd566_1 CB@8_mAd566_2 CB@8_mAd567_1 
+CB@8_mAd567_2 CB@8_mAd570_1 CB@8_mAd570_2 CB@8_mAd571_1 CB@8_mAd571_2 CB@8_mAd572_1 CB@8_mAd572_2 CB@8_mAd573_1 CB@8_mAd573_2 CB@8_mAd575_1 CB@8_mAd575_2 CB@8_mAd576_1 CB@8_mAd576_2 CB@8_mAd577_1 CB@8_mAd577_2 CB@8_mAd600_1 CB@8_mAd600_2 CB@8_mAd601_1 CB@8_mAd601_2 CB@8_mAd602_1 CB@8_mAd602_2 CB@8_mAd604_1 CB@8_mAd604_2 CB@8_mAd605_1 CB@8_mAd605_2 CB@8_mAd606_1 CB@8_mAd606_2 CB@8_mAd607_1 CB@8_mAd607_2 CB@8_mAd610_1 CB@8_mAd610_2 CB@8_mAd611_1 CB@8_mAd611_2 CB@8_mAd612_1 CB@8_mAd612_2 CB@8_mAd613_1 
+CB@8_mAd613_2 CB@8_mAd614_1 CB@8_mAd614_2 CB@8_mAd615_1 CB@8_mAd615_2 CB@8_mAd616_1 CB@8_mAd616_2 CB@8_mAd617_1 CB@8_mAd617_2 CB@8_mAd620_1 CB@8_mAd620_2 CB@8_mAd621_1 CB@8_mAd621_2 CB@8_mAd622_1 CB@8_mAd622_2 CB@8_mAd623_1 CB@8_mAd623_2 CB@8_mAd624_1 CB@8_mAd624_2 CB@8_mAd625_1 CB@8_mAd625_2 CB@8_mAd626_1 CB@8_mAd626_2 CB@8_mAd627_1 CB@8_mAd627_2 CB@8_mAd630_1 CB@8_mAd630_2 CB@8_mAd631_1 CB@8_mAd631_2 CB@8_mAd632_1 CB@8_mAd632_2 CB@8_mAd633_1 CB@8_mAd633_2 CB@8_mAd634_1 CB@8_mAd634_2 CB@8_mAd635_1 
+CB@8_mAd635_2 CB@8_mAd636_1 CB@8_mAd636_2 CB@8_mAd637_1 CB@8_mAd637_2 CB@8_mAd640_1 CB@8_mAd640_2 CB@8_mAd641_1 CB@8_mAd641_2 CB@8_mAd642_1 CB@8_mAd642_2 CB@8_mAd643_1 CB@8_mAd643_2 CB@8_mAd644_1 CB@8_mAd644_2 CB@8_mAd645_1 CB@8_mAd645_2 CB@8_mAd646_1 CB@8_mAd646_2 CB@8_mAd647_1 CB@8_mAd647_2 CB@8_mAd650_1 CB@8_mAd650_2 CB@8_mAd651_1 CB@8_mAd651_2 CB@8_mAd652_1 CB@8_mAd652_2 CB@8_mAd653_1 CB@8_mAd653_2 CB@8_mAd654_1 CB@8_mAd654_2 CB@8_mAd655_1 CB@8_mAd655_2 CB@8_mAd656_1 CB@8_mAd656_2 CB@8_mAd657_1 
+CB@8_mAd657_2 CB@8_mAd660_1 CB@8_mAd660_2 CB@8_mAd661_1 CB@8_mAd661_2 CB@8_mAd662_1 CB@8_mAd662_2 CB@8_mAd663_1 CB@8_mAd663_2 CB@8_mAd664_1 CB@8_mAd664_2 CB@8_mAd665_1 CB@8_mAd665_2 CB@8_mAd666_1 CB@8_mAd666_2 CB@8_mAd667_1 CB@8_mAd667_2 CB@8_mAd675_1 CB@8_mAd675_2 CB@8_mAd676_1 CB@8_mAd676_2 CB@8_mAd677_1 CB@8_mAd677_2 CB@8_mAd700_1 CB@8_mAd700_2 CB@8_mAd710_1 CB@8_mAd710_2 CB@8_mAd711_1 CB@8_mAd711_2 CB@8_mAd717_1 CB@8_mAd717_2 CB@8_mAd720_1 CB@8_mAd720_2 CB@8_mAd721_1 CB@8_mAd721_2 CB@8_mAd722_1 
+CB@8_mAd722_2 CB@8_mAd723_1 CB@8_mAd723_2 CB@8_mAd724_1 CB@8_mAd724_2 CB@8_mAd725_1 CB@8_mAd725_2 CB@8_mAd726_1 CB@8_mAd726_2 CB@8_mAd727_1 CB@8_mAd727_2 CB@8_mAd730_1 CB@8_mAd730_2 CB@8_mAd731_1 CB@8_mAd731_2 CB@8_mAd732_1 CB@8_mAd732_2 CB@8_mAd733_1 CB@8_mAd733_2 CB@8_mAd734_1 CB@8_mAd734_2 CB@8_mAd735_1 CB@8_mAd735_2 CB@8_mAd736_1 CB@8_mAd736_2 CB@8_mAd737_1 CB@8_mAd737_2 CB@8_mAd740_1 CB@8_mAd740_2 CB@8_mAd741_1 CB@8_mAd741_2 CB@8_mAd742_1 CB@8_mAd742_2 CB@8_mAd743_1 CB@8_mAd743_2 CB@8_mAd744_1 
+CB@8_mAd744_2 CB@8_mAd745_1 CB@8_mAd745_2 CB@8_mAd746_1 CB@8_mAd746_2 CB@8_mAd747_1 CB@8_mAd747_2 CB@8_mAd750_1 CB@8_mAd750_2 CB@8_mAd751_1 CB@8_mAd751_2 CB@8_mAd752_1 CB@8_mAd752_2 CB@8_mAd753_1 CB@8_mAd753_2 CB@8_mAd754_1 CB@8_mAd754_2 CB@8_mAd755_1 CB@8_mAd755_2 CB@8_mAd756_1 CB@8_mAd756_2 CB@8_mAd757_1 CB@8_mAd757_2 CB@8_mAd760_1 CB@8_mAd760_2 CB@8_mAd761_1 CB@8_mAd761_2 CB@8_mAd762_1 CB@8_mAd762_2 CB@8_mAd763_1 CB@8_mAd763_2 CB@8_mAd764_1 CB@8_mAd764_2 CB@8_mAd765_1 CB@8_mAd765_2 CB@8_mAd766_1 
+CB@8_mAd766_2 CB@8_mAd767_1 CB@8_mAd767_2 CB@8_mAd771_1 CB@8_mAd771_2 CB@8_mAd772_1 CB@8_mAd772_2 CB@8_mAd773_1 CB@8_mAd773_2 CB@8_mAd774_1 CB@8_mAd774_2 CB@8_mAd775_1 CB@8_mAd775_2 CB@8_mAd776_1 CB@8_mAd776_2 CB@8_mAd777_1 CB@8_mAd777_2 CB@8_X0 CB@8_X1 CB@8_X10 CB@8_X11 CB@8_X12 CB@8_X13 CB@8_X2 CB@8_X3 CB@8_X4 CB@8_X5 CB@8_X6 CB@8_X7 CB@8_X8 CB@8_X9 CB@8_Y1 CB@8_Y10 CB@8_Y11 CB@8_Y12 CB@8_Y2 CB@8_Y3 CB@8_Y4 CB@8_Y5 CB@8_Y6 CB@8_Y7 CB@8_Y8 CB@8_Y9 CB@8_Z1 CB@8_Z10 CB@8_Z11 CB@8_Z12 CB@8_Z2 CB@8_Z3 CB@8_Z4 
+CB@8_Z5 CB@8_Z6 CB@8_Z7 CB@8_Z8 CB@8_Z9 _5400TP094__CB
XCB@9 CB@9_K0 CB@9_K1 CB@9_K10 CB@9_K11 CB@9_K12 CB@9_K13 CB@9_K2 CB@9_K3 CB@9_K4 CB@9_K5 CB@9_K6 CB@9_K7 CB@9_K8 CB@9_K9 CB@9_mAd000_1 CB@9_mAd000_2 CB@9_mAd001_1 CB@9_mAd001_2 CB@9_mAd002_1 CB@9_mAd002_2 CB@9_mAd003_1 CB@9_mAd003_2 CB@9_mAd004_1 CB@9_mAd004_2 CB@9_mAd005_1 CB@9_mAd005_2 CB@9_mAd006_1 CB@9_mAd006_2 CB@9_mAd007_1 CB@9_mAd007_2 CB@9_mAd010_1 CB@9_mAd010_2 CB@9_mAd011_1 CB@9_mAd011_2 CB@9_mAd012_1 CB@9_mAd012_2 CB@9_mAd013_1 CB@9_mAd013_2 CB@9_mAd014_1 CB@9_mAd014_2 CB@9_mAd015_1 
+CB@9_mAd015_2 CB@9_mAd016_1 CB@9_mAd016_2 CB@9_mAd017_1 CB@9_mAd017_2 CB@9_mAd020_1 CB@9_mAd020_2 CB@9_mAd021_1 CB@9_mAd021_2 CB@9_mAd022_1 CB@9_mAd022_2 CB@9_mAd023_1 CB@9_mAd023_2 CB@9_mAd024_1 CB@9_mAd024_2 CB@9_mAd025_1 CB@9_mAd025_2 CB@9_mAd026_1 CB@9_mAd026_2 CB@9_mAd027_1 CB@9_mAd027_2 CB@9_mAd030_1 CB@9_mAd030_2 CB@9_mAd031_1 CB@9_mAd031_2 CB@9_mAd032_1 CB@9_mAd032_2 CB@9_mAd033_1 CB@9_mAd033_2 CB@9_mAd034_1 CB@9_mAd034_2 CB@9_mAd035_1 CB@9_mAd035_2 CB@9_mAd036_1 CB@9_mAd036_2 CB@9_mAd037_1 
+CB@9_mAd037_2 CB@9_mAd040_1 CB@9_mAd040_2 CB@9_mAd041_1 CB@9_mAd041_2 CB@9_mAd042_1 CB@9_mAd042_2 CB@9_mAd043_1 CB@9_mAd043_2 CB@9_mAd044_1 CB@9_mAd044_2 CB@9_mAd045_1 CB@9_mAd045_2 CB@9_mAd046_1 CB@9_mAd046_2 CB@9_mAd047_1 CB@9_mAd047_2 CB@9_mAd050_1 CB@9_mAd050_2 CB@9_mAd051_1 CB@9_mAd051_2 CB@9_mAd052_1 CB@9_mAd052_2 CB@9_mAd053_1 CB@9_mAd053_2 CB@9_mAd054_1 CB@9_mAd054_2 CB@9_mAd055_1 CB@9_mAd055_2 CB@9_mAd056_1 CB@9_mAd056_2 CB@9_mAd057_1 CB@9_mAd057_2 CB@9_mAd060_1 CB@9_mAd060_2 CB@9_mAd066_1 
+CB@9_mAd066_2 CB@9_mAd067_1 CB@9_mAd067_2 CB@9_mAd100_1 CB@9_mAd100_2 CB@9_mAd101_1 CB@9_mAd101_2 CB@9_mAd102_1 CB@9_mAd102_2 CB@9_mAd110_1 CB@9_mAd110_2 CB@9_mAd111_1 CB@9_mAd111_2 CB@9_mAd112_1 CB@9_mAd112_2 CB@9_mAd113_1 CB@9_mAd113_2 CB@9_mAd114_1 CB@9_mAd114_2 CB@9_mAd115_1 CB@9_mAd115_2 CB@9_mAd116_1 CB@9_mAd116_2 CB@9_mAd117_1 CB@9_mAd117_2 CB@9_mAd120_1 CB@9_mAd120_2 CB@9_mAd121_1 CB@9_mAd121_2 CB@9_mAd122_1 CB@9_mAd122_2 CB@9_mAd123_1 CB@9_mAd123_2 CB@9_mAd124_1 CB@9_mAd124_2 CB@9_mAd125_1 
+CB@9_mAd125_2 CB@9_mAd126_1 CB@9_mAd126_2 CB@9_mAd127_1 CB@9_mAd127_2 CB@9_mAd130_1 CB@9_mAd130_2 CB@9_mAd131_1 CB@9_mAd131_2 CB@9_mAd132_1 CB@9_mAd132_2 CB@9_mAd133_1 CB@9_mAd133_2 CB@9_mAd134_1 CB@9_mAd134_2 CB@9_mAd135_1 CB@9_mAd135_2 CB@9_mAd136_1 CB@9_mAd136_2 CB@9_mAd137_1 CB@9_mAd137_2 CB@9_mAd140_1 CB@9_mAd140_2 CB@9_mAd141_1 CB@9_mAd141_2 CB@9_mAd142_1 CB@9_mAd142_2 CB@9_mAd143_1 CB@9_mAd143_2 CB@9_mAd144_1 CB@9_mAd144_2 CB@9_mAd145_1 CB@9_mAd145_2 CB@9_mAd146_1 CB@9_mAd146_2 CB@9_mAd147_1 
+CB@9_mAd147_2 CB@9_mAd150_1 CB@9_mAd150_2 CB@9_mAd151_1 CB@9_mAd151_2 CB@9_mAd152_1 CB@9_mAd152_2 CB@9_mAd153_1 CB@9_mAd153_2 CB@9_mAd154_1 CB@9_mAd154_2 CB@9_mAd155_1 CB@9_mAd155_2 CB@9_mAd156_1 CB@9_mAd156_2 CB@9_mAd157_1 CB@9_mAd157_2 CB@9_mAd160_1 CB@9_mAd160_2 CB@9_mAd161_1 CB@9_mAd161_2 CB@9_mAd162_1 CB@9_mAd162_2 CB@9_mAd163_1 CB@9_mAd163_2 CB@9_mAd164_1 CB@9_mAd164_2 CB@9_mAd165_1 CB@9_mAd165_2 CB@9_mAd166_1 CB@9_mAd166_2 CB@9_mAd167_1 CB@9_mAd167_2 CB@9_mAd170_1 CB@9_mAd170_2 CB@9_mAd171_1 
+CB@9_mAd171_2 CB@9_mAd172_1 CB@9_mAd172_2 CB@9_mAd173_1 CB@9_mAd173_2 CB@9_mAd175_1 CB@9_mAd175_2 CB@9_mAd176_1 CB@9_mAd176_2 CB@9_mAd177_1 CB@9_mAd177_2 CB@9_mAd200_1 CB@9_mAd200_2 CB@9_mAd201_1 CB@9_mAd201_2 CB@9_mAd202_1 CB@9_mAd202_2 CB@9_mAd204_1 CB@9_mAd204_2 CB@9_mAd205_1 CB@9_mAd205_2 CB@9_mAd206_1 CB@9_mAd206_2 CB@9_mAd207_1 CB@9_mAd207_2 CB@9_mAd210_1 CB@9_mAd210_2 CB@9_mAd211_1 CB@9_mAd211_2 CB@9_mAd212_1 CB@9_mAd212_2 CB@9_mAd213_1 CB@9_mAd213_2 CB@9_mAd214_1 CB@9_mAd214_2 CB@9_mAd215_1 
+CB@9_mAd215_2 CB@9_mAd216_1 CB@9_mAd216_2 CB@9_mAd217_1 CB@9_mAd217_2 CB@9_mAd220_1 CB@9_mAd220_2 CB@9_mAd221_1 CB@9_mAd221_2 CB@9_mAd222_1 CB@9_mAd222_2 CB@9_mAd223_1 CB@9_mAd223_2 CB@9_mAd224_1 CB@9_mAd224_2 CB@9_mAd225_1 CB@9_mAd225_2 CB@9_mAd226_1 CB@9_mAd226_2 CB@9_mAd227_1 CB@9_mAd227_2 CB@9_mAd230_1 CB@9_mAd230_2 CB@9_mAd231_1 CB@9_mAd231_2 CB@9_mAd232_1 CB@9_mAd232_2 CB@9_mAd233_1 CB@9_mAd233_2 CB@9_mAd234_1 CB@9_mAd234_2 CB@9_mAd235_1 CB@9_mAd235_2 CB@9_mAd236_1 CB@9_mAd236_2 CB@9_mAd237_1 
+CB@9_mAd237_2 CB@9_mAd240_1 CB@9_mAd240_2 CB@9_mAd241_1 CB@9_mAd241_2 CB@9_mAd242_1 CB@9_mAd242_2 CB@9_mAd243_1 CB@9_mAd243_2 CB@9_mAd244_1 CB@9_mAd244_2 CB@9_mAd245_1 CB@9_mAd245_2 CB@9_mAd246_1 CB@9_mAd246_2 CB@9_mAd247_1 CB@9_mAd247_2 CB@9_mAd250_1 CB@9_mAd250_2 CB@9_mAd251_1 CB@9_mAd251_2 CB@9_mAd252_1 CB@9_mAd252_2 CB@9_mAd253_1 CB@9_mAd253_2 CB@9_mAd254_1 CB@9_mAd254_2 CB@9_mAd255_1 CB@9_mAd255_2 CB@9_mAd256_1 CB@9_mAd256_2 CB@9_mAd257_1 CB@9_mAd257_2 CB@9_mAd260_1 CB@9_mAd260_2 CB@9_mAd261_1 
+CB@9_mAd261_2 CB@9_mAd262_1 CB@9_mAd262_2 CB@9_mAd263_1 CB@9_mAd263_2 CB@9_mAd264_1 CB@9_mAd264_2 CB@9_mAd265_1 CB@9_mAd265_2 CB@9_mAd266_1 CB@9_mAd266_2 CB@9_mAd267_1 CB@9_mAd267_2 CB@9_mAd275_1 CB@9_mAd275_2 CB@9_mAd276_1 CB@9_mAd276_2 CB@9_mAd277_1 CB@9_mAd277_2 CB@9_mAd300_1 CB@9_mAd300_2 CB@9_mAd310_1 CB@9_mAd310_2 CB@9_mAd311_1 CB@9_mAd311_2 CB@9_mAd317_1 CB@9_mAd317_2 CB@9_mAd320_1 CB@9_mAd320_2 CB@9_mAd321_1 CB@9_mAd321_2 CB@9_mAd322_1 CB@9_mAd322_2 CB@9_mAd323_1 CB@9_mAd323_2 CB@9_mAd324_1 
+CB@9_mAd324_2 CB@9_mAd325_1 CB@9_mAd325_2 CB@9_mAd326_1 CB@9_mAd326_2 CB@9_mAd327_1 CB@9_mAd327_2 CB@9_mAd330_1 CB@9_mAd330_2 CB@9_mAd331_1 CB@9_mAd331_2 CB@9_mAd332_1 CB@9_mAd332_2 CB@9_mAd333_1 CB@9_mAd333_2 CB@9_mAd334_1 CB@9_mAd334_2 CB@9_mAd335_1 CB@9_mAd335_2 CB@9_mAd336_1 CB@9_mAd336_2 CB@9_mAd337_1 CB@9_mAd337_2 CB@9_mAd340_1 CB@9_mAd340_2 CB@9_mAd341_1 CB@9_mAd341_2 CB@9_mAd342_1 CB@9_mAd342_2 CB@9_mAd343_1 CB@9_mAd343_2 CB@9_mAd344_1 CB@9_mAd344_2 CB@9_mAd345_1 CB@9_mAd345_2 CB@9_mAd346_1 
+CB@9_mAd346_2 CB@9_mAd347_1 CB@9_mAd347_2 CB@9_mAd350_1 CB@9_mAd350_2 CB@9_mAd351_1 CB@9_mAd351_2 CB@9_mAd352_1 CB@9_mAd352_2 CB@9_mAd353_1 CB@9_mAd353_2 CB@9_mAd354_1 CB@9_mAd354_2 CB@9_mAd355_1 CB@9_mAd355_2 CB@9_mAd356_1 CB@9_mAd356_2 CB@9_mAd357_1 CB@9_mAd357_2 CB@9_mAd360_1 CB@9_mAd360_2 CB@9_mAd361_1 CB@9_mAd361_2 CB@9_mAd362_1 CB@9_mAd362_2 CB@9_mAd363_1 CB@9_mAd363_2 CB@9_mAd364_1 CB@9_mAd364_2 CB@9_mAd365_1 CB@9_mAd365_2 CB@9_mAd366_1 CB@9_mAd366_2 CB@9_mAd367_1 CB@9_mAd367_2 CB@9_mAd371_1 
+CB@9_mAd371_2 CB@9_mAd372_1 CB@9_mAd372_2 CB@9_mAd373_1 CB@9_mAd373_2 CB@9_mAd374_1 CB@9_mAd374_2 CB@9_mAd375_1 CB@9_mAd375_2 CB@9_mAd376_1 CB@9_mAd376_2 CB@9_mAd377_1 CB@9_mAd377_2 CB@9_mAd400_1 CB@9_mAd400_2 CB@9_mAd401_1 CB@9_mAd401_2 CB@9_mAd402_1 CB@9_mAd402_2 CB@9_mAd403_1 CB@9_mAd403_2 CB@9_mAd404_1 CB@9_mAd404_2 CB@9_mAd405_1 CB@9_mAd405_2 CB@9_mAd406_1 CB@9_mAd406_2 CB@9_mAd407_1 CB@9_mAd407_2 CB@9_mAd410_1 CB@9_mAd410_2 CB@9_mAd411_1 CB@9_mAd411_2 CB@9_mAd412_1 CB@9_mAd412_2 CB@9_mAd413_1 
+CB@9_mAd413_2 CB@9_mAd414_1 CB@9_mAd414_2 CB@9_mAd415_1 CB@9_mAd415_2 CB@9_mAd416_1 CB@9_mAd416_2 CB@9_mAd417_1 CB@9_mAd417_2 CB@9_mAd420_1 CB@9_mAd420_2 CB@9_mAd421_1 CB@9_mAd421_2 CB@9_mAd422_1 CB@9_mAd422_2 CB@9_mAd423_1 CB@9_mAd423_2 CB@9_mAd424_1 CB@9_mAd424_2 CB@9_mAd425_1 CB@9_mAd425_2 CB@9_mAd426_1 CB@9_mAd426_2 CB@9_mAd427_1 CB@9_mAd427_2 CB@9_mAd430_1 CB@9_mAd430_2 CB@9_mAd431_1 CB@9_mAd431_2 CB@9_mAd432_1 CB@9_mAd432_2 CB@9_mAd433_1 CB@9_mAd433_2 CB@9_mAd434_1 CB@9_mAd434_2 CB@9_mAd435_1 
+CB@9_mAd435_2 CB@9_mAd436_1 CB@9_mAd436_2 CB@9_mAd437_1 CB@9_mAd437_2 CB@9_mAd440_1 CB@9_mAd440_2 CB@9_mAd441_1 CB@9_mAd441_2 CB@9_mAd442_1 CB@9_mAd442_2 CB@9_mAd443_1 CB@9_mAd443_2 CB@9_mAd444_1 CB@9_mAd444_2 CB@9_mAd445_1 CB@9_mAd445_2 CB@9_mAd446_1 CB@9_mAd446_2 CB@9_mAd447_1 CB@9_mAd447_2 CB@9_mAd450_1 CB@9_mAd450_2 CB@9_mAd451_1 CB@9_mAd451_2 CB@9_mAd452_1 CB@9_mAd452_2 CB@9_mAd453_1 CB@9_mAd453_2 CB@9_mAd454_1 CB@9_mAd454_2 CB@9_mAd455_1 CB@9_mAd455_2 CB@9_mAd456_1 CB@9_mAd456_2 CB@9_mAd457_1 
+CB@9_mAd457_2 CB@9_mAd460_1 CB@9_mAd460_2 CB@9_mAd466_1 CB@9_mAd466_2 CB@9_mAd467_1 CB@9_mAd467_2 CB@9_mAd500_1 CB@9_mAd500_2 CB@9_mAd501_1 CB@9_mAd501_2 CB@9_mAd502_1 CB@9_mAd502_2 CB@9_mAd508_1 CB@9_mAd508_2 CB@9_mAd509_1 CB@9_mAd509_2 CB@9_mAd512_1 CB@9_mAd512_2 CB@9_mAd513_1 CB@9_mAd513_2 CB@9_mAd514_1 CB@9_mAd514_2 CB@9_mAd515_1 CB@9_mAd515_2 CB@9_mAd516_1 CB@9_mAd516_2 CB@9_mAd517_1 CB@9_mAd517_2 CB@9_mAd520_1 CB@9_mAd520_2 CB@9_mAd521_1 CB@9_mAd521_2 CB@9_mAd522_1 CB@9_mAd522_2 CB@9_mAd523_1 
+CB@9_mAd523_2 CB@9_mAd524_1 CB@9_mAd524_2 CB@9_mAd525_1 CB@9_mAd525_2 CB@9_mAd526_1 CB@9_mAd526_2 CB@9_mAd527_1 CB@9_mAd527_2 CB@9_mAd530_1 CB@9_mAd530_2 CB@9_mAd531_1 CB@9_mAd531_2 CB@9_mAd532_1 CB@9_mAd532_2 CB@9_mAd533_1 CB@9_mAd533_2 CB@9_mAd534_1 CB@9_mAd534_2 CB@9_mAd535_1 CB@9_mAd535_2 CB@9_mAd536_1 CB@9_mAd536_2 CB@9_mAd537_1 CB@9_mAd537_2 CB@9_mAd540_1 CB@9_mAd540_2 CB@9_mAd541_1 CB@9_mAd541_2 CB@9_mAd542_1 CB@9_mAd542_2 CB@9_mAd543_1 CB@9_mAd543_2 CB@9_mAd544_1 CB@9_mAd544_2 CB@9_mAd545_1 
+CB@9_mAd545_2 CB@9_mAd546_1 CB@9_mAd546_2 CB@9_mAd547_1 CB@9_mAd547_2 CB@9_mAd550_1 CB@9_mAd550_2 CB@9_mAd551_1 CB@9_mAd551_2 CB@9_mAd552_1 CB@9_mAd552_2 CB@9_mAd553_1 CB@9_mAd553_2 CB@9_mAd554_1 CB@9_mAd554_2 CB@9_mAd555_1 CB@9_mAd555_2 CB@9_mAd556_1 CB@9_mAd556_2 CB@9_mAd557_1 CB@9_mAd557_2 CB@9_mAd560_1 CB@9_mAd560_2 CB@9_mAd561_1 CB@9_mAd561_2 CB@9_mAd562_1 CB@9_mAd562_2 CB@9_mAd563_1 CB@9_mAd563_2 CB@9_mAd564_1 CB@9_mAd564_2 CB@9_mAd565_1 CB@9_mAd565_2 CB@9_mAd566_1 CB@9_mAd566_2 CB@9_mAd567_1 
+CB@9_mAd567_2 CB@9_mAd570_1 CB@9_mAd570_2 CB@9_mAd571_1 CB@9_mAd571_2 CB@9_mAd572_1 CB@9_mAd572_2 CB@9_mAd573_1 CB@9_mAd573_2 CB@9_mAd575_1 CB@9_mAd575_2 CB@9_mAd576_1 CB@9_mAd576_2 CB@9_mAd577_1 CB@9_mAd577_2 CB@9_mAd600_1 CB@9_mAd600_2 CB@9_mAd601_1 CB@9_mAd601_2 CB@9_mAd602_1 CB@9_mAd602_2 CB@9_mAd604_1 CB@9_mAd604_2 CB@9_mAd605_1 CB@9_mAd605_2 CB@9_mAd606_1 CB@9_mAd606_2 CB@9_mAd607_1 CB@9_mAd607_2 CB@9_mAd610_1 CB@9_mAd610_2 CB@9_mAd611_1 CB@9_mAd611_2 CB@9_mAd612_1 CB@9_mAd612_2 CB@9_mAd613_1 
+CB@9_mAd613_2 CB@9_mAd614_1 CB@9_mAd614_2 CB@9_mAd615_1 CB@9_mAd615_2 CB@9_mAd616_1 CB@9_mAd616_2 CB@9_mAd617_1 CB@9_mAd617_2 CB@9_mAd620_1 CB@9_mAd620_2 CB@9_mAd621_1 CB@9_mAd621_2 CB@9_mAd622_1 CB@9_mAd622_2 CB@9_mAd623_1 CB@9_mAd623_2 CB@9_mAd624_1 CB@9_mAd624_2 CB@9_mAd625_1 CB@9_mAd625_2 CB@9_mAd626_1 CB@9_mAd626_2 CB@9_mAd627_1 CB@9_mAd627_2 CB@9_mAd630_1 CB@9_mAd630_2 CB@9_mAd631_1 CB@9_mAd631_2 CB@9_mAd632_1 CB@9_mAd632_2 CB@9_mAd633_1 CB@9_mAd633_2 CB@9_mAd634_1 CB@9_mAd634_2 CB@9_mAd635_1 
+CB@9_mAd635_2 CB@9_mAd636_1 CB@9_mAd636_2 CB@9_mAd637_1 CB@9_mAd637_2 CB@9_mAd640_1 CB@9_mAd640_2 CB@9_mAd641_1 CB@9_mAd641_2 CB@9_mAd642_1 CB@9_mAd642_2 CB@9_mAd643_1 CB@9_mAd643_2 CB@9_mAd644_1 CB@9_mAd644_2 CB@9_mAd645_1 CB@9_mAd645_2 CB@9_mAd646_1 CB@9_mAd646_2 CB@9_mAd647_1 CB@9_mAd647_2 CB@9_mAd650_1 CB@9_mAd650_2 CB@9_mAd651_1 CB@9_mAd651_2 CB@9_mAd652_1 CB@9_mAd652_2 CB@9_mAd653_1 CB@9_mAd653_2 CB@9_mAd654_1 CB@9_mAd654_2 CB@9_mAd655_1 CB@9_mAd655_2 CB@9_mAd656_1 CB@9_mAd656_2 CB@9_mAd657_1 
+CB@9_mAd657_2 CB@9_mAd660_1 CB@9_mAd660_2 CB@9_mAd661_1 CB@9_mAd661_2 CB@9_mAd662_1 CB@9_mAd662_2 CB@9_mAd663_1 CB@9_mAd663_2 CB@9_mAd664_1 CB@9_mAd664_2 CB@9_mAd665_1 CB@9_mAd665_2 CB@9_mAd666_1 CB@9_mAd666_2 CB@9_mAd667_1 CB@9_mAd667_2 CB@9_mAd675_1 CB@9_mAd675_2 CB@9_mAd676_1 CB@9_mAd676_2 CB@9_mAd677_1 CB@9_mAd677_2 CB@9_mAd700_1 CB@9_mAd700_2 CB@9_mAd710_1 CB@9_mAd710_2 CB@9_mAd711_1 CB@9_mAd711_2 CB@9_mAd717_1 CB@9_mAd717_2 CB@9_mAd720_1 CB@9_mAd720_2 CB@9_mAd721_1 CB@9_mAd721_2 CB@9_mAd722_1 
+CB@9_mAd722_2 CB@9_mAd723_1 CB@9_mAd723_2 CB@9_mAd724_1 CB@9_mAd724_2 CB@9_mAd725_1 CB@9_mAd725_2 CB@9_mAd726_1 CB@9_mAd726_2 CB@9_mAd727_1 CB@9_mAd727_2 CB@9_mAd730_1 CB@9_mAd730_2 CB@9_mAd731_1 CB@9_mAd731_2 CB@9_mAd732_1 CB@9_mAd732_2 CB@9_mAd733_1 CB@9_mAd733_2 CB@9_mAd734_1 CB@9_mAd734_2 CB@9_mAd735_1 CB@9_mAd735_2 CB@9_mAd736_1 CB@9_mAd736_2 CB@9_mAd737_1 CB@9_mAd737_2 CB@9_mAd740_1 CB@9_mAd740_2 CB@9_mAd741_1 CB@9_mAd741_2 CB@9_mAd742_1 CB@9_mAd742_2 CB@9_mAd743_1 CB@9_mAd743_2 CB@9_mAd744_1 
+CB@9_mAd744_2 CB@9_mAd745_1 CB@9_mAd745_2 CB@9_mAd746_1 CB@9_mAd746_2 CB@9_mAd747_1 CB@9_mAd747_2 CB@9_mAd750_1 CB@9_mAd750_2 CB@9_mAd751_1 CB@9_mAd751_2 CB@9_mAd752_1 CB@9_mAd752_2 CB@9_mAd753_1 CB@9_mAd753_2 CB@9_mAd754_1 CB@9_mAd754_2 CB@9_mAd755_1 CB@9_mAd755_2 CB@9_mAd756_1 CB@9_mAd756_2 CB@9_mAd757_1 CB@9_mAd757_2 CB@9_mAd760_1 CB@9_mAd760_2 CB@9_mAd761_1 CB@9_mAd761_2 CB@9_mAd762_1 CB@9_mAd762_2 CB@9_mAd763_1 CB@9_mAd763_2 CB@9_mAd764_1 CB@9_mAd764_2 CB@9_mAd765_1 CB@9_mAd765_2 CB@9_mAd766_1 
+CB@9_mAd766_2 CB@9_mAd767_1 CB@9_mAd767_2 CB@9_mAd771_1 CB@9_mAd771_2 CB@9_mAd772_1 CB@9_mAd772_2 CB@9_mAd773_1 CB@9_mAd773_2 CB@9_mAd774_1 CB@9_mAd774_2 CB@9_mAd775_1 CB@9_mAd775_2 CB@9_mAd776_1 CB@9_mAd776_2 CB@9_mAd777_1 CB@9_mAd777_2 CB@9_X0 CB@9_X1 CB@9_X10 CB@9_X11 CB@9_X12 CB@9_X13 CB@9_X2 CB@9_X3 CB@9_X4 CB@9_X5 CB@9_X6 CB@9_X7 CB@9_X8 CB@9_X9 CB@9_Y1 CB@9_Y10 CB@9_Y11 CB@9_Y12 CB@9_Y2 CB@9_Y3 CB@9_Y4 CB@9_Y5 CB@9_Y6 CB@9_Y7 CB@9_Y8 CB@9_Y9 CB@9_Z1 CB@9_Z10 CB@9_Z11 CB@9_Z12 CB@9_Z2 CB@9_Z3 CB@9_Z4 
+CB@9_Z5 CB@9_Z6 CB@9_Z7 CB@9_Z8 CB@9_Z9 _5400TP094__CB
XCB@10 CB@10_K0 CB@10_K1 CB@10_K10 CB@10_K11 CB@10_K12 CB@10_K13 CB@10_K2 CB@10_K3 CB@10_K4 CB@10_K5 CB@10_K6 CB@10_K7 CB@10_K8 CB@10_K9 CB@10_mAd000_1 CB@10_mAd000_2 CB@10_mAd001_1 CB@10_mAd001_2 CB@10_mAd002_1 CB@10_mAd002_2 CB@10_mAd003_1 CB@10_mAd003_2 CB@10_mAd004_1 CB@10_mAd004_2 CB@10_mAd005_1 CB@10_mAd005_2 CB@10_mAd006_1 CB@10_mAd006_2 CB@10_mAd007_1 CB@10_mAd007_2 CB@10_mAd010_1 CB@10_mAd010_2 CB@10_mAd011_1 CB@10_mAd011_2 CB@10_mAd012_1 CB@10_mAd012_2 CB@10_mAd013_1 CB@10_mAd013_2 CB@10_mAd014_1 
+CB@10_mAd014_2 CB@10_mAd015_1 CB@10_mAd015_2 CB@10_mAd016_1 CB@10_mAd016_2 CB@10_mAd017_1 CB@10_mAd017_2 CB@10_mAd020_1 CB@10_mAd020_2 CB@10_mAd021_1 CB@10_mAd021_2 CB@10_mAd022_1 CB@10_mAd022_2 CB@10_mAd023_1 CB@10_mAd023_2 CB@10_mAd024_1 CB@10_mAd024_2 CB@10_mAd025_1 CB@10_mAd025_2 CB@10_mAd026_1 CB@10_mAd026_2 CB@10_mAd027_1 CB@10_mAd027_2 CB@10_mAd030_1 CB@10_mAd030_2 CB@10_mAd031_1 CB@10_mAd031_2 CB@10_mAd032_1 CB@10_mAd032_2 CB@10_mAd033_1 CB@10_mAd033_2 CB@10_mAd034_1 CB@10_mAd034_2 CB@10_mAd035_1 
+CB@10_mAd035_2 CB@10_mAd036_1 CB@10_mAd036_2 CB@10_mAd037_1 CB@10_mAd037_2 CB@10_mAd040_1 CB@10_mAd040_2 CB@10_mAd041_1 CB@10_mAd041_2 CB@10_mAd042_1 CB@10_mAd042_2 CB@10_mAd043_1 CB@10_mAd043_2 CB@10_mAd044_1 CB@10_mAd044_2 CB@10_mAd045_1 CB@10_mAd045_2 CB@10_mAd046_1 CB@10_mAd046_2 CB@10_mAd047_1 CB@10_mAd047_2 CB@10_mAd050_1 CB@10_mAd050_2 CB@10_mAd051_1 CB@10_mAd051_2 CB@10_mAd052_1 CB@10_mAd052_2 CB@10_mAd053_1 CB@10_mAd053_2 CB@10_mAd054_1 CB@10_mAd054_2 CB@10_mAd055_1 CB@10_mAd055_2 CB@10_mAd056_1 
+CB@10_mAd056_2 CB@10_mAd057_1 CB@10_mAd057_2 CB@10_mAd060_1 CB@10_mAd060_2 CB@10_mAd066_1 CB@10_mAd066_2 CB@10_mAd067_1 CB@10_mAd067_2 CB@10_mAd100_1 CB@10_mAd100_2 CB@10_mAd101_1 CB@10_mAd101_2 CB@10_mAd102_1 CB@10_mAd102_2 CB@10_mAd110_1 CB@10_mAd110_2 CB@10_mAd111_1 CB@10_mAd111_2 CB@10_mAd112_1 CB@10_mAd112_2 CB@10_mAd113_1 CB@10_mAd113_2 CB@10_mAd114_1 CB@10_mAd114_2 CB@10_mAd115_1 CB@10_mAd115_2 CB@10_mAd116_1 CB@10_mAd116_2 CB@10_mAd117_1 CB@10_mAd117_2 CB@10_mAd120_1 CB@10_mAd120_2 CB@10_mAd121_1 
+CB@10_mAd121_2 CB@10_mAd122_1 CB@10_mAd122_2 CB@10_mAd123_1 CB@10_mAd123_2 CB@10_mAd124_1 CB@10_mAd124_2 CB@10_mAd125_1 CB@10_mAd125_2 CB@10_mAd126_1 CB@10_mAd126_2 CB@10_mAd127_1 CB@10_mAd127_2 CB@10_mAd130_1 CB@10_mAd130_2 CB@10_mAd131_1 CB@10_mAd131_2 CB@10_mAd132_1 CB@10_mAd132_2 CB@10_mAd133_1 CB@10_mAd133_2 CB@10_mAd134_1 CB@10_mAd134_2 CB@10_mAd135_1 CB@10_mAd135_2 CB@10_mAd136_1 CB@10_mAd136_2 CB@10_mAd137_1 CB@10_mAd137_2 CB@10_mAd140_1 CB@10_mAd140_2 CB@10_mAd141_1 CB@10_mAd141_2 CB@10_mAd142_1 
+CB@10_mAd142_2 CB@10_mAd143_1 CB@10_mAd143_2 CB@10_mAd144_1 CB@10_mAd144_2 CB@10_mAd145_1 CB@10_mAd145_2 CB@10_mAd146_1 CB@10_mAd146_2 CB@10_mAd147_1 CB@10_mAd147_2 CB@10_mAd150_1 CB@10_mAd150_2 CB@10_mAd151_1 CB@10_mAd151_2 CB@10_mAd152_1 CB@10_mAd152_2 CB@10_mAd153_1 CB@10_mAd153_2 CB@10_mAd154_1 CB@10_mAd154_2 CB@10_mAd155_1 CB@10_mAd155_2 CB@10_mAd156_1 CB@10_mAd156_2 CB@10_mAd157_1 CB@10_mAd157_2 CB@10_mAd160_1 CB@10_mAd160_2 CB@10_mAd161_1 CB@10_mAd161_2 CB@10_mAd162_1 CB@10_mAd162_2 CB@10_mAd163_1 
+CB@10_mAd163_2 CB@10_mAd164_1 CB@10_mAd164_2 CB@10_mAd165_1 CB@10_mAd165_2 CB@10_mAd166_1 CB@10_mAd166_2 CB@10_mAd167_1 CB@10_mAd167_2 CB@10_mAd170_1 CB@10_mAd170_2 CB@10_mAd171_1 CB@10_mAd171_2 CB@10_mAd172_1 CB@10_mAd172_2 CB@10_mAd173_1 CB@10_mAd173_2 CB@10_mAd175_1 CB@10_mAd175_2 CB@10_mAd176_1 CB@10_mAd176_2 CB@10_mAd177_1 CB@10_mAd177_2 CB@10_mAd200_1 CB@10_mAd200_2 CB@10_mAd201_1 CB@10_mAd201_2 CB@10_mAd202_1 CB@10_mAd202_2 CB@10_mAd204_1 CB@10_mAd204_2 CB@10_mAd205_1 CB@10_mAd205_2 CB@10_mAd206_1 
+CB@10_mAd206_2 CB@10_mAd207_1 CB@10_mAd207_2 CB@10_mAd210_1 CB@10_mAd210_2 CB@10_mAd211_1 CB@10_mAd211_2 CB@10_mAd212_1 CB@10_mAd212_2 CB@10_mAd213_1 CB@10_mAd213_2 CB@10_mAd214_1 CB@10_mAd214_2 CB@10_mAd215_1 CB@10_mAd215_2 CB@10_mAd216_1 CB@10_mAd216_2 CB@10_mAd217_1 CB@10_mAd217_2 CB@10_mAd220_1 CB@10_mAd220_2 CB@10_mAd221_1 CB@10_mAd221_2 CB@10_mAd222_1 CB@10_mAd222_2 CB@10_mAd223_1 CB@10_mAd223_2 CB@10_mAd224_1 CB@10_mAd224_2 CB@10_mAd225_1 CB@10_mAd225_2 CB@10_mAd226_1 CB@10_mAd226_2 CB@10_mAd227_1 
+CB@10_mAd227_2 CB@10_mAd230_1 CB@10_mAd230_2 CB@10_mAd231_1 CB@10_mAd231_2 CB@10_mAd232_1 CB@10_mAd232_2 CB@10_mAd233_1 CB@10_mAd233_2 CB@10_mAd234_1 CB@10_mAd234_2 CB@10_mAd235_1 CB@10_mAd235_2 CB@10_mAd236_1 CB@10_mAd236_2 CB@10_mAd237_1 CB@10_mAd237_2 CB@10_mAd240_1 CB@10_mAd240_2 CB@10_mAd241_1 CB@10_mAd241_2 CB@10_mAd242_1 CB@10_mAd242_2 CB@10_mAd243_1 CB@10_mAd243_2 CB@10_mAd244_1 CB@10_mAd244_2 CB@10_mAd245_1 CB@10_mAd245_2 CB@10_mAd246_1 CB@10_mAd246_2 CB@10_mAd247_1 CB@10_mAd247_2 CB@10_mAd250_1 
+CB@10_mAd250_2 CB@10_mAd251_1 CB@10_mAd251_2 CB@10_mAd252_1 CB@10_mAd252_2 CB@10_mAd253_1 CB@10_mAd253_2 CB@10_mAd254_1 CB@10_mAd254_2 CB@10_mAd255_1 CB@10_mAd255_2 CB@10_mAd256_1 CB@10_mAd256_2 CB@10_mAd257_1 CB@10_mAd257_2 CB@10_mAd260_1 CB@10_mAd260_2 CB@10_mAd261_1 CB@10_mAd261_2 CB@10_mAd262_1 CB@10_mAd262_2 CB@10_mAd263_1 CB@10_mAd263_2 CB@10_mAd264_1 CB@10_mAd264_2 CB@10_mAd265_1 CB@10_mAd265_2 CB@10_mAd266_1 CB@10_mAd266_2 CB@10_mAd267_1 CB@10_mAd267_2 CB@10_mAd275_1 CB@10_mAd275_2 CB@10_mAd276_1 
+CB@10_mAd276_2 CB@10_mAd277_1 CB@10_mAd277_2 CB@10_mAd300_1 CB@10_mAd300_2 CB@10_mAd310_1 CB@10_mAd310_2 CB@10_mAd311_1 CB@10_mAd311_2 CB@10_mAd317_1 CB@10_mAd317_2 CB@10_mAd320_1 CB@10_mAd320_2 CB@10_mAd321_1 CB@10_mAd321_2 CB@10_mAd322_1 CB@10_mAd322_2 CB@10_mAd323_1 CB@10_mAd323_2 CB@10_mAd324_1 CB@10_mAd324_2 CB@10_mAd325_1 CB@10_mAd325_2 CB@10_mAd326_1 CB@10_mAd326_2 CB@10_mAd327_1 CB@10_mAd327_2 CB@10_mAd330_1 CB@10_mAd330_2 CB@10_mAd331_1 CB@10_mAd331_2 CB@10_mAd332_1 CB@10_mAd332_2 CB@10_mAd333_1 
+CB@10_mAd333_2 CB@10_mAd334_1 CB@10_mAd334_2 CB@10_mAd335_1 CB@10_mAd335_2 CB@10_mAd336_1 CB@10_mAd336_2 CB@10_mAd337_1 CB@10_mAd337_2 CB@10_mAd340_1 CB@10_mAd340_2 CB@10_mAd341_1 CB@10_mAd341_2 CB@10_mAd342_1 CB@10_mAd342_2 CB@10_mAd343_1 CB@10_mAd343_2 CB@10_mAd344_1 CB@10_mAd344_2 CB@10_mAd345_1 CB@10_mAd345_2 CB@10_mAd346_1 CB@10_mAd346_2 CB@10_mAd347_1 CB@10_mAd347_2 CB@10_mAd350_1 CB@10_mAd350_2 CB@10_mAd351_1 CB@10_mAd351_2 CB@10_mAd352_1 CB@10_mAd352_2 CB@10_mAd353_1 CB@10_mAd353_2 CB@10_mAd354_1 
+CB@10_mAd354_2 CB@10_mAd355_1 CB@10_mAd355_2 CB@10_mAd356_1 CB@10_mAd356_2 CB@10_mAd357_1 CB@10_mAd357_2 CB@10_mAd360_1 CB@10_mAd360_2 CB@10_mAd361_1 CB@10_mAd361_2 CB@10_mAd362_1 CB@10_mAd362_2 CB@10_mAd363_1 CB@10_mAd363_2 CB@10_mAd364_1 CB@10_mAd364_2 CB@10_mAd365_1 CB@10_mAd365_2 CB@10_mAd366_1 CB@10_mAd366_2 CB@10_mAd367_1 CB@10_mAd367_2 CB@10_mAd371_1 CB@10_mAd371_2 CB@10_mAd372_1 CB@10_mAd372_2 CB@10_mAd373_1 CB@10_mAd373_2 CB@10_mAd374_1 CB@10_mAd374_2 CB@10_mAd375_1 CB@10_mAd375_2 CB@10_mAd376_1 
+CB@10_mAd376_2 CB@10_mAd377_1 CB@10_mAd377_2 CB@10_mAd400_1 CB@10_mAd400_2 CB@10_mAd401_1 CB@10_mAd401_2 CB@10_mAd402_1 CB@10_mAd402_2 CB@10_mAd403_1 CB@10_mAd403_2 CB@10_mAd404_1 CB@10_mAd404_2 CB@10_mAd405_1 CB@10_mAd405_2 CB@10_mAd406_1 CB@10_mAd406_2 CB@10_mAd407_1 CB@10_mAd407_2 CB@10_mAd410_1 CB@10_mAd410_2 CB@10_mAd411_1 CB@10_mAd411_2 CB@10_mAd412_1 CB@10_mAd412_2 CB@10_mAd413_1 CB@10_mAd413_2 CB@10_mAd414_1 CB@10_mAd414_2 CB@10_mAd415_1 CB@10_mAd415_2 CB@10_mAd416_1 CB@10_mAd416_2 CB@10_mAd417_1 
+CB@10_mAd417_2 CB@10_mAd420_1 CB@10_mAd420_2 CB@10_mAd421_1 CB@10_mAd421_2 CB@10_mAd422_1 CB@10_mAd422_2 CB@10_mAd423_1 CB@10_mAd423_2 CB@10_mAd424_1 CB@10_mAd424_2 CB@10_mAd425_1 CB@10_mAd425_2 CB@10_mAd426_1 CB@10_mAd426_2 CB@10_mAd427_1 CB@10_mAd427_2 CB@10_mAd430_1 CB@10_mAd430_2 CB@10_mAd431_1 CB@10_mAd431_2 CB@10_mAd432_1 CB@10_mAd432_2 CB@10_mAd433_1 CB@10_mAd433_2 CB@10_mAd434_1 CB@10_mAd434_2 CB@10_mAd435_1 CB@10_mAd435_2 CB@10_mAd436_1 CB@10_mAd436_2 CB@10_mAd437_1 CB@10_mAd437_2 CB@10_mAd440_1 
+CB@10_mAd440_2 CB@10_mAd441_1 CB@10_mAd441_2 CB@10_mAd442_1 CB@10_mAd442_2 CB@10_mAd443_1 CB@10_mAd443_2 CB@10_mAd444_1 CB@10_mAd444_2 CB@10_mAd445_1 CB@10_mAd445_2 CB@10_mAd446_1 CB@10_mAd446_2 CB@10_mAd447_1 CB@10_mAd447_2 CB@10_mAd450_1 CB@10_mAd450_2 CB@10_mAd451_1 CB@10_mAd451_2 CB@10_mAd452_1 CB@10_mAd452_2 CB@10_mAd453_1 CB@10_mAd453_2 CB@10_mAd454_1 CB@10_mAd454_2 CB@10_mAd455_1 CB@10_mAd455_2 CB@10_mAd456_1 CB@10_mAd456_2 CB@10_mAd457_1 CB@10_mAd457_2 CB@10_mAd460_1 CB@10_mAd460_2 CB@10_mAd466_1 
+CB@10_mAd466_2 CB@10_mAd467_1 CB@10_mAd467_2 CB@10_mAd500_1 CB@10_mAd500_2 CB@10_mAd501_1 CB@10_mAd501_2 CB@10_mAd502_1 CB@10_mAd502_2 CB@10_mAd508_1 CB@10_mAd508_2 CB@10_mAd509_1 CB@10_mAd509_2 CB@10_mAd512_1 CB@10_mAd512_2 CB@10_mAd513_1 CB@10_mAd513_2 CB@10_mAd514_1 CB@10_mAd514_2 CB@10_mAd515_1 CB@10_mAd515_2 CB@10_mAd516_1 CB@10_mAd516_2 CB@10_mAd517_1 CB@10_mAd517_2 CB@10_mAd520_1 CB@10_mAd520_2 CB@10_mAd521_1 CB@10_mAd521_2 CB@10_mAd522_1 CB@10_mAd522_2 CB@10_mAd523_1 CB@10_mAd523_2 CB@10_mAd524_1 
+CB@10_mAd524_2 CB@10_mAd525_1 CB@10_mAd525_2 CB@10_mAd526_1 CB@10_mAd526_2 CB@10_mAd527_1 CB@10_mAd527_2 CB@10_mAd530_1 CB@10_mAd530_2 CB@10_mAd531_1 CB@10_mAd531_2 CB@10_mAd532_1 CB@10_mAd532_2 CB@10_mAd533_1 CB@10_mAd533_2 CB@10_mAd534_1 CB@10_mAd534_2 CB@10_mAd535_1 CB@10_mAd535_2 CB@10_mAd536_1 CB@10_mAd536_2 CB@10_mAd537_1 CB@10_mAd537_2 CB@10_mAd540_1 CB@10_mAd540_2 CB@10_mAd541_1 CB@10_mAd541_2 CB@10_mAd542_1 CB@10_mAd542_2 CB@10_mAd543_1 CB@10_mAd543_2 CB@10_mAd544_1 CB@10_mAd544_2 CB@10_mAd545_1 
+CB@10_mAd545_2 CB@10_mAd546_1 CB@10_mAd546_2 CB@10_mAd547_1 CB@10_mAd547_2 CB@10_mAd550_1 CB@10_mAd550_2 CB@10_mAd551_1 CB@10_mAd551_2 CB@10_mAd552_1 CB@10_mAd552_2 CB@10_mAd553_1 CB@10_mAd553_2 CB@10_mAd554_1 CB@10_mAd554_2 CB@10_mAd555_1 CB@10_mAd555_2 CB@10_mAd556_1 CB@10_mAd556_2 CB@10_mAd557_1 CB@10_mAd557_2 CB@10_mAd560_1 CB@10_mAd560_2 CB@10_mAd561_1 CB@10_mAd561_2 CB@10_mAd562_1 CB@10_mAd562_2 CB@10_mAd563_1 CB@10_mAd563_2 CB@10_mAd564_1 CB@10_mAd564_2 CB@10_mAd565_1 CB@10_mAd565_2 CB@10_mAd566_1 
+CB@10_mAd566_2 CB@10_mAd567_1 CB@10_mAd567_2 CB@10_mAd570_1 CB@10_mAd570_2 CB@10_mAd571_1 CB@10_mAd571_2 CB@10_mAd572_1 CB@10_mAd572_2 CB@10_mAd573_1 CB@10_mAd573_2 CB@10_mAd575_1 CB@10_mAd575_2 CB@10_mAd576_1 CB@10_mAd576_2 CB@10_mAd577_1 CB@10_mAd577_2 CB@10_mAd600_1 CB@10_mAd600_2 CB@10_mAd601_1 CB@10_mAd601_2 CB@10_mAd602_1 CB@10_mAd602_2 CB@10_mAd604_1 CB@10_mAd604_2 CB@10_mAd605_1 CB@10_mAd605_2 CB@10_mAd606_1 CB@10_mAd606_2 CB@10_mAd607_1 CB@10_mAd607_2 CB@10_mAd610_1 CB@10_mAd610_2 CB@10_mAd611_1 
+CB@10_mAd611_2 CB@10_mAd612_1 CB@10_mAd612_2 CB@10_mAd613_1 CB@10_mAd613_2 CB@10_mAd614_1 CB@10_mAd614_2 CB@10_mAd615_1 CB@10_mAd615_2 CB@10_mAd616_1 CB@10_mAd616_2 CB@10_mAd617_1 CB@10_mAd617_2 CB@10_mAd620_1 CB@10_mAd620_2 CB@10_mAd621_1 CB@10_mAd621_2 CB@10_mAd622_1 CB@10_mAd622_2 CB@10_mAd623_1 CB@10_mAd623_2 CB@10_mAd624_1 CB@10_mAd624_2 CB@10_mAd625_1 CB@10_mAd625_2 CB@10_mAd626_1 CB@10_mAd626_2 CB@10_mAd627_1 CB@10_mAd627_2 CB@10_mAd630_1 CB@10_mAd630_2 CB@10_mAd631_1 CB@10_mAd631_2 CB@10_mAd632_1 
+CB@10_mAd632_2 CB@10_mAd633_1 CB@10_mAd633_2 CB@10_mAd634_1 CB@10_mAd634_2 CB@10_mAd635_1 CB@10_mAd635_2 CB@10_mAd636_1 CB@10_mAd636_2 CB@10_mAd637_1 CB@10_mAd637_2 CB@10_mAd640_1 CB@10_mAd640_2 CB@10_mAd641_1 CB@10_mAd641_2 CB@10_mAd642_1 CB@10_mAd642_2 CB@10_mAd643_1 CB@10_mAd643_2 CB@10_mAd644_1 CB@10_mAd644_2 CB@10_mAd645_1 CB@10_mAd645_2 CB@10_mAd646_1 CB@10_mAd646_2 CB@10_mAd647_1 CB@10_mAd647_2 CB@10_mAd650_1 CB@10_mAd650_2 CB@10_mAd651_1 CB@10_mAd651_2 CB@10_mAd652_1 CB@10_mAd652_2 CB@10_mAd653_1 
+CB@10_mAd653_2 CB@10_mAd654_1 CB@10_mAd654_2 CB@10_mAd655_1 CB@10_mAd655_2 CB@10_mAd656_1 CB@10_mAd656_2 CB@10_mAd657_1 CB@10_mAd657_2 CB@10_mAd660_1 CB@10_mAd660_2 CB@10_mAd661_1 CB@10_mAd661_2 CB@10_mAd662_1 CB@10_mAd662_2 CB@10_mAd663_1 CB@10_mAd663_2 CB@10_mAd664_1 CB@10_mAd664_2 CB@10_mAd665_1 CB@10_mAd665_2 CB@10_mAd666_1 CB@10_mAd666_2 CB@10_mAd667_1 CB@10_mAd667_2 CB@10_mAd675_1 CB@10_mAd675_2 CB@10_mAd676_1 CB@10_mAd676_2 CB@10_mAd677_1 CB@10_mAd677_2 CB@10_mAd700_1 CB@10_mAd700_2 CB@10_mAd710_1 
+CB@10_mAd710_2 CB@10_mAd711_1 CB@10_mAd711_2 CB@10_mAd717_1 CB@10_mAd717_2 CB@10_mAd720_1 CB@10_mAd720_2 CB@10_mAd721_1 CB@10_mAd721_2 CB@10_mAd722_1 CB@10_mAd722_2 CB@10_mAd723_1 CB@10_mAd723_2 CB@10_mAd724_1 CB@10_mAd724_2 CB@10_mAd725_1 CB@10_mAd725_2 CB@10_mAd726_1 CB@10_mAd726_2 CB@10_mAd727_1 CB@10_mAd727_2 CB@10_mAd730_1 CB@10_mAd730_2 CB@10_mAd731_1 CB@10_mAd731_2 CB@10_mAd732_1 CB@10_mAd732_2 CB@10_mAd733_1 CB@10_mAd733_2 CB@10_mAd734_1 CB@10_mAd734_2 CB@10_mAd735_1 CB@10_mAd735_2 CB@10_mAd736_1 
+CB@10_mAd736_2 CB@10_mAd737_1 CB@10_mAd737_2 CB@10_mAd740_1 CB@10_mAd740_2 CB@10_mAd741_1 CB@10_mAd741_2 CB@10_mAd742_1 CB@10_mAd742_2 CB@10_mAd743_1 CB@10_mAd743_2 CB@10_mAd744_1 CB@10_mAd744_2 CB@10_mAd745_1 CB@10_mAd745_2 CB@10_mAd746_1 CB@10_mAd746_2 CB@10_mAd747_1 CB@10_mAd747_2 CB@10_mAd750_1 CB@10_mAd750_2 CB@10_mAd751_1 CB@10_mAd751_2 CB@10_mAd752_1 CB@10_mAd752_2 CB@10_mAd753_1 CB@10_mAd753_2 CB@10_mAd754_1 CB@10_mAd754_2 CB@10_mAd755_1 CB@10_mAd755_2 CB@10_mAd756_1 CB@10_mAd756_2 CB@10_mAd757_1 
+CB@10_mAd757_2 CB@10_mAd760_1 CB@10_mAd760_2 CB@10_mAd761_1 CB@10_mAd761_2 CB@10_mAd762_1 CB@10_mAd762_2 CB@10_mAd763_1 CB@10_mAd763_2 CB@10_mAd764_1 CB@10_mAd764_2 CB@10_mAd765_1 CB@10_mAd765_2 CB@10_mAd766_1 CB@10_mAd766_2 CB@10_mAd767_1 CB@10_mAd767_2 CB@10_mAd771_1 CB@10_mAd771_2 CB@10_mAd772_1 CB@10_mAd772_2 CB@10_mAd773_1 CB@10_mAd773_2 CB@10_mAd774_1 CB@10_mAd774_2 CB@10_mAd775_1 CB@10_mAd775_2 CB@10_mAd776_1 CB@10_mAd776_2 CB@10_mAd777_1 CB@10_mAd777_2 CB@10_X0 CB@10_X1 CB@10_X10 CB@10_X11 
+CB@10_X12 CB@10_X13 CB@10_X2 CB@10_X3 CB@10_X4 CB@10_X5 CB@10_X6 CB@10_X7 CB@10_X8 CB@10_X9 CB@10_Y1 CB@10_Y10 CB@10_Y11 CB@10_Y12 CB@10_Y2 CB@10_Y3 CB@10_Y4 CB@10_Y5 CB@10_Y6 CB@10_Y7 CB@10_Y8 CB@10_Y9 CB@10_Z1 CB@10_Z10 CB@10_Z11 CB@10_Z12 CB@10_Z2 CB@10_Z3 CB@10_Z4 CB@10_Z5 CB@10_Z6 CB@10_Z7 CB@10_Z8 CB@10_Z9 _5400TP094__CB
XCB@11 CB@11_K0 CB@11_K1 CB@11_K10 CB@11_K11 CB@11_K12 CB@11_K13 CB@11_K2 CB@11_K3 CB@11_K4 CB@11_K5 CB@11_K6 CB@11_K7 CB@11_K8 CB@11_K9 CB@11_mAd000_1 CB@11_mAd000_2 CB@11_mAd001_1 CB@11_mAd001_2 CB@11_mAd002_1 CB@11_mAd002_2 CB@11_mAd003_1 CB@11_mAd003_2 CB@11_mAd004_1 CB@11_mAd004_2 CB@11_mAd005_1 CB@11_mAd005_2 CB@11_mAd006_1 CB@11_mAd006_2 CB@11_mAd007_1 CB@11_mAd007_2 CB@11_mAd010_1 CB@11_mAd010_2 CB@11_mAd011_1 CB@11_mAd011_2 CB@11_mAd012_1 CB@11_mAd012_2 CB@11_mAd013_1 CB@11_mAd013_2 CB@11_mAd014_1 
+CB@11_mAd014_2 CB@11_mAd015_1 CB@11_mAd015_2 CB@11_mAd016_1 CB@11_mAd016_2 CB@11_mAd017_1 CB@11_mAd017_2 CB@11_mAd020_1 CB@11_mAd020_2 CB@11_mAd021_1 CB@11_mAd021_2 CB@11_mAd022_1 CB@11_mAd022_2 CB@11_mAd023_1 CB@11_mAd023_2 CB@11_mAd024_1 CB@11_mAd024_2 CB@11_mAd025_1 CB@11_mAd025_2 CB@11_mAd026_1 CB@11_mAd026_2 CB@11_mAd027_1 CB@11_mAd027_2 CB@11_mAd030_1 CB@11_mAd030_2 CB@11_mAd031_1 CB@11_mAd031_2 CB@11_mAd032_1 CB@11_mAd032_2 CB@11_mAd033_1 CB@11_mAd033_2 CB@11_mAd034_1 CB@11_mAd034_2 CB@11_mAd035_1 
+CB@11_mAd035_2 CB@11_mAd036_1 CB@11_mAd036_2 CB@11_mAd037_1 CB@11_mAd037_2 CB@11_mAd040_1 CB@11_mAd040_2 CB@11_mAd041_1 CB@11_mAd041_2 CB@11_mAd042_1 CB@11_mAd042_2 CB@11_mAd043_1 CB@11_mAd043_2 CB@11_mAd044_1 CB@11_mAd044_2 CB@11_mAd045_1 CB@11_mAd045_2 CB@11_mAd046_1 CB@11_mAd046_2 CB@11_mAd047_1 CB@11_mAd047_2 CB@11_mAd050_1 CB@11_mAd050_2 CB@11_mAd051_1 CB@11_mAd051_2 CB@11_mAd052_1 CB@11_mAd052_2 CB@11_mAd053_1 CB@11_mAd053_2 CB@11_mAd054_1 CB@11_mAd054_2 CB@11_mAd055_1 CB@11_mAd055_2 CB@11_mAd056_1 
+CB@11_mAd056_2 CB@11_mAd057_1 CB@11_mAd057_2 CB@11_mAd060_1 CB@11_mAd060_2 CB@11_mAd066_1 CB@11_mAd066_2 CB@11_mAd067_1 CB@11_mAd067_2 CB@11_mAd100_1 CB@11_mAd100_2 CB@11_mAd101_1 CB@11_mAd101_2 CB@11_mAd102_1 CB@11_mAd102_2 CB@11_mAd110_1 CB@11_mAd110_2 CB@11_mAd111_1 CB@11_mAd111_2 CB@11_mAd112_1 CB@11_mAd112_2 CB@11_mAd113_1 CB@11_mAd113_2 CB@11_mAd114_1 CB@11_mAd114_2 CB@11_mAd115_1 CB@11_mAd115_2 CB@11_mAd116_1 CB@11_mAd116_2 CB@11_mAd117_1 CB@11_mAd117_2 CB@11_mAd120_1 CB@11_mAd120_2 CB@11_mAd121_1 
+CB@11_mAd121_2 CB@11_mAd122_1 CB@11_mAd122_2 CB@11_mAd123_1 CB@11_mAd123_2 CB@11_mAd124_1 CB@11_mAd124_2 CB@11_mAd125_1 CB@11_mAd125_2 CB@11_mAd126_1 CB@11_mAd126_2 CB@11_mAd127_1 CB@11_mAd127_2 CB@11_mAd130_1 CB@11_mAd130_2 CB@11_mAd131_1 CB@11_mAd131_2 CB@11_mAd132_1 CB@11_mAd132_2 CB@11_mAd133_1 CB@11_mAd133_2 CB@11_mAd134_1 CB@11_mAd134_2 CB@11_mAd135_1 CB@11_mAd135_2 CB@11_mAd136_1 CB@11_mAd136_2 CB@11_mAd137_1 CB@11_mAd137_2 CB@11_mAd140_1 CB@11_mAd140_2 CB@11_mAd141_1 CB@11_mAd141_2 CB@11_mAd142_1 
+CB@11_mAd142_2 CB@11_mAd143_1 CB@11_mAd143_2 CB@11_mAd144_1 CB@11_mAd144_2 CB@11_mAd145_1 CB@11_mAd145_2 CB@11_mAd146_1 CB@11_mAd146_2 CB@11_mAd147_1 CB@11_mAd147_2 CB@11_mAd150_1 CB@11_mAd150_2 CB@11_mAd151_1 CB@11_mAd151_2 CB@11_mAd152_1 CB@11_mAd152_2 CB@11_mAd153_1 CB@11_mAd153_2 CB@11_mAd154_1 CB@11_mAd154_2 CB@11_mAd155_1 CB@11_mAd155_2 CB@11_mAd156_1 CB@11_mAd156_2 CB@11_mAd157_1 CB@11_mAd157_2 CB@11_mAd160_1 CB@11_mAd160_2 CB@11_mAd161_1 CB@11_mAd161_2 CB@11_mAd162_1 CB@11_mAd162_2 CB@11_mAd163_1 
+CB@11_mAd163_2 CB@11_mAd164_1 CB@11_mAd164_2 CB@11_mAd165_1 CB@11_mAd165_2 CB@11_mAd166_1 CB@11_mAd166_2 CB@11_mAd167_1 CB@11_mAd167_2 CB@11_mAd170_1 CB@11_mAd170_2 CB@11_mAd171_1 CB@11_mAd171_2 CB@11_mAd172_1 CB@11_mAd172_2 CB@11_mAd173_1 CB@11_mAd173_2 CB@11_mAd175_1 CB@11_mAd175_2 CB@11_mAd176_1 CB@11_mAd176_2 CB@11_mAd177_1 CB@11_mAd177_2 CB@11_mAd200_1 CB@11_mAd200_2 CB@11_mAd201_1 CB@11_mAd201_2 CB@11_mAd202_1 CB@11_mAd202_2 CB@11_mAd204_1 CB@11_mAd204_2 CB@11_mAd205_1 CB@11_mAd205_2 CB@11_mAd206_1 
+CB@11_mAd206_2 CB@11_mAd207_1 CB@11_mAd207_2 CB@11_mAd210_1 CB@11_mAd210_2 CB@11_mAd211_1 CB@11_mAd211_2 CB@11_mAd212_1 CB@11_mAd212_2 CB@11_mAd213_1 CB@11_mAd213_2 CB@11_mAd214_1 CB@11_mAd214_2 CB@11_mAd215_1 CB@11_mAd215_2 CB@11_mAd216_1 CB@11_mAd216_2 CB@11_mAd217_1 CB@11_mAd217_2 CB@11_mAd220_1 CB@11_mAd220_2 CB@11_mAd221_1 CB@11_mAd221_2 CB@11_mAd222_1 CB@11_mAd222_2 CB@11_mAd223_1 CB@11_mAd223_2 CB@11_mAd224_1 CB@11_mAd224_2 CB@11_mAd225_1 CB@11_mAd225_2 CB@11_mAd226_1 CB@11_mAd226_2 CB@11_mAd227_1 
+CB@11_mAd227_2 CB@11_mAd230_1 CB@11_mAd230_2 CB@11_mAd231_1 CB@11_mAd231_2 CB@11_mAd232_1 CB@11_mAd232_2 CB@11_mAd233_1 CB@11_mAd233_2 CB@11_mAd234_1 CB@11_mAd234_2 CB@11_mAd235_1 CB@11_mAd235_2 CB@11_mAd236_1 CB@11_mAd236_2 CB@11_mAd237_1 CB@11_mAd237_2 CB@11_mAd240_1 CB@11_mAd240_2 CB@11_mAd241_1 CB@11_mAd241_2 CB@11_mAd242_1 CB@11_mAd242_2 CB@11_mAd243_1 CB@11_mAd243_2 CB@11_mAd244_1 CB@11_mAd244_2 CB@11_mAd245_1 CB@11_mAd245_2 CB@11_mAd246_1 CB@11_mAd246_2 CB@11_mAd247_1 CB@11_mAd247_2 CB@11_mAd250_1 
+CB@11_mAd250_2 CB@11_mAd251_1 CB@11_mAd251_2 CB@11_mAd252_1 CB@11_mAd252_2 CB@11_mAd253_1 CB@11_mAd253_2 CB@11_mAd254_1 CB@11_mAd254_2 CB@11_mAd255_1 CB@11_mAd255_2 CB@11_mAd256_1 CB@11_mAd256_2 CB@11_mAd257_1 CB@11_mAd257_2 CB@11_mAd260_1 CB@11_mAd260_2 CB@11_mAd261_1 CB@11_mAd261_2 CB@11_mAd262_1 CB@11_mAd262_2 CB@11_mAd263_1 CB@11_mAd263_2 CB@11_mAd264_1 CB@11_mAd264_2 CB@11_mAd265_1 CB@11_mAd265_2 CB@11_mAd266_1 CB@11_mAd266_2 CB@11_mAd267_1 CB@11_mAd267_2 CB@11_mAd275_1 CB@11_mAd275_2 CB@11_mAd276_1 
+CB@11_mAd276_2 CB@11_mAd277_1 CB@11_mAd277_2 CB@11_mAd300_1 CB@11_mAd300_2 CB@11_mAd310_1 CB@11_mAd310_2 CB@11_mAd311_1 CB@11_mAd311_2 CB@11_mAd317_1 CB@11_mAd317_2 CB@11_mAd320_1 CB@11_mAd320_2 CB@11_mAd321_1 CB@11_mAd321_2 CB@11_mAd322_1 CB@11_mAd322_2 CB@11_mAd323_1 CB@11_mAd323_2 CB@11_mAd324_1 CB@11_mAd324_2 CB@11_mAd325_1 CB@11_mAd325_2 CB@11_mAd326_1 CB@11_mAd326_2 CB@11_mAd327_1 CB@11_mAd327_2 CB@11_mAd330_1 CB@11_mAd330_2 CB@11_mAd331_1 CB@11_mAd331_2 CB@11_mAd332_1 CB@11_mAd332_2 CB@11_mAd333_1 
+CB@11_mAd333_2 CB@11_mAd334_1 CB@11_mAd334_2 CB@11_mAd335_1 CB@11_mAd335_2 CB@11_mAd336_1 CB@11_mAd336_2 CB@11_mAd337_1 CB@11_mAd337_2 CB@11_mAd340_1 CB@11_mAd340_2 CB@11_mAd341_1 CB@11_mAd341_2 CB@11_mAd342_1 CB@11_mAd342_2 CB@11_mAd343_1 CB@11_mAd343_2 CB@11_mAd344_1 CB@11_mAd344_2 CB@11_mAd345_1 CB@11_mAd345_2 CB@11_mAd346_1 CB@11_mAd346_2 CB@11_mAd347_1 CB@11_mAd347_2 CB@11_mAd350_1 CB@11_mAd350_2 CB@11_mAd351_1 CB@11_mAd351_2 CB@11_mAd352_1 CB@11_mAd352_2 CB@11_mAd353_1 CB@11_mAd353_2 CB@11_mAd354_1 
+CB@11_mAd354_2 CB@11_mAd355_1 CB@11_mAd355_2 CB@11_mAd356_1 CB@11_mAd356_2 CB@11_mAd357_1 CB@11_mAd357_2 CB@11_mAd360_1 CB@11_mAd360_2 CB@11_mAd361_1 CB@11_mAd361_2 CB@11_mAd362_1 CB@11_mAd362_2 CB@11_mAd363_1 CB@11_mAd363_2 CB@11_mAd364_1 CB@11_mAd364_2 CB@11_mAd365_1 CB@11_mAd365_2 CB@11_mAd366_1 CB@11_mAd366_2 CB@11_mAd367_1 CB@11_mAd367_2 CB@11_mAd371_1 CB@11_mAd371_2 CB@11_mAd372_1 CB@11_mAd372_2 CB@11_mAd373_1 CB@11_mAd373_2 CB@11_mAd374_1 CB@11_mAd374_2 CB@11_mAd375_1 CB@11_mAd375_2 CB@11_mAd376_1 
+CB@11_mAd376_2 CB@11_mAd377_1 CB@11_mAd377_2 CB@11_mAd400_1 CB@11_mAd400_2 CB@11_mAd401_1 CB@11_mAd401_2 CB@11_mAd402_1 CB@11_mAd402_2 CB@11_mAd403_1 CB@11_mAd403_2 CB@11_mAd404_1 CB@11_mAd404_2 CB@11_mAd405_1 CB@11_mAd405_2 CB@11_mAd406_1 CB@11_mAd406_2 CB@11_mAd407_1 CB@11_mAd407_2 CB@11_mAd410_1 CB@11_mAd410_2 CB@11_mAd411_1 CB@11_mAd411_2 CB@11_mAd412_1 CB@11_mAd412_2 CB@11_mAd413_1 CB@11_mAd413_2 CB@11_mAd414_1 CB@11_mAd414_2 CB@11_mAd415_1 CB@11_mAd415_2 CB@11_mAd416_1 CB@11_mAd416_2 CB@11_mAd417_1 
+CB@11_mAd417_2 CB@11_mAd420_1 CB@11_mAd420_2 CB@11_mAd421_1 CB@11_mAd421_2 CB@11_mAd422_1 CB@11_mAd422_2 CB@11_mAd423_1 CB@11_mAd423_2 CB@11_mAd424_1 CB@11_mAd424_2 CB@11_mAd425_1 CB@11_mAd425_2 CB@11_mAd426_1 CB@11_mAd426_2 CB@11_mAd427_1 CB@11_mAd427_2 CB@11_mAd430_1 CB@11_mAd430_2 CB@11_mAd431_1 CB@11_mAd431_2 CB@11_mAd432_1 CB@11_mAd432_2 CB@11_mAd433_1 CB@11_mAd433_2 CB@11_mAd434_1 CB@11_mAd434_2 CB@11_mAd435_1 CB@11_mAd435_2 CB@11_mAd436_1 CB@11_mAd436_2 CB@11_mAd437_1 CB@11_mAd437_2 CB@11_mAd440_1 
+CB@11_mAd440_2 CB@11_mAd441_1 CB@11_mAd441_2 CB@11_mAd442_1 CB@11_mAd442_2 CB@11_mAd443_1 CB@11_mAd443_2 CB@11_mAd444_1 CB@11_mAd444_2 CB@11_mAd445_1 CB@11_mAd445_2 CB@11_mAd446_1 CB@11_mAd446_2 CB@11_mAd447_1 CB@11_mAd447_2 CB@11_mAd450_1 CB@11_mAd450_2 CB@11_mAd451_1 CB@11_mAd451_2 CB@11_mAd452_1 CB@11_mAd452_2 CB@11_mAd453_1 CB@11_mAd453_2 CB@11_mAd454_1 CB@11_mAd454_2 CB@11_mAd455_1 CB@11_mAd455_2 CB@11_mAd456_1 CB@11_mAd456_2 CB@11_mAd457_1 CB@11_mAd457_2 CB@11_mAd460_1 CB@11_mAd460_2 CB@11_mAd466_1 
+CB@11_mAd466_2 CB@11_mAd467_1 CB@11_mAd467_2 CB@11_mAd500_1 CB@11_mAd500_2 CB@11_mAd501_1 CB@11_mAd501_2 CB@11_mAd502_1 CB@11_mAd502_2 CB@11_mAd508_1 CB@11_mAd508_2 CB@11_mAd509_1 CB@11_mAd509_2 CB@11_mAd512_1 CB@11_mAd512_2 CB@11_mAd513_1 CB@11_mAd513_2 CB@11_mAd514_1 CB@11_mAd514_2 CB@11_mAd515_1 CB@11_mAd515_2 CB@11_mAd516_1 CB@11_mAd516_2 CB@11_mAd517_1 CB@11_mAd517_2 CB@11_mAd520_1 CB@11_mAd520_2 CB@11_mAd521_1 CB@11_mAd521_2 CB@11_mAd522_1 CB@11_mAd522_2 CB@11_mAd523_1 CB@11_mAd523_2 CB@11_mAd524_1 
+CB@11_mAd524_2 CB@11_mAd525_1 CB@11_mAd525_2 CB@11_mAd526_1 CB@11_mAd526_2 CB@11_mAd527_1 CB@11_mAd527_2 CB@11_mAd530_1 CB@11_mAd530_2 CB@11_mAd531_1 CB@11_mAd531_2 CB@11_mAd532_1 CB@11_mAd532_2 CB@11_mAd533_1 CB@11_mAd533_2 CB@11_mAd534_1 CB@11_mAd534_2 CB@11_mAd535_1 CB@11_mAd535_2 CB@11_mAd536_1 CB@11_mAd536_2 CB@11_mAd537_1 CB@11_mAd537_2 CB@11_mAd540_1 CB@11_mAd540_2 CB@11_mAd541_1 CB@11_mAd541_2 CB@11_mAd542_1 CB@11_mAd542_2 CB@11_mAd543_1 CB@11_mAd543_2 CB@11_mAd544_1 CB@11_mAd544_2 CB@11_mAd545_1 
+CB@11_mAd545_2 CB@11_mAd546_1 CB@11_mAd546_2 CB@11_mAd547_1 CB@11_mAd547_2 CB@11_mAd550_1 CB@11_mAd550_2 CB@11_mAd551_1 CB@11_mAd551_2 CB@11_mAd552_1 CB@11_mAd552_2 CB@11_mAd553_1 CB@11_mAd553_2 CB@11_mAd554_1 CB@11_mAd554_2 CB@11_mAd555_1 CB@11_mAd555_2 CB@11_mAd556_1 CB@11_mAd556_2 CB@11_mAd557_1 CB@11_mAd557_2 CB@11_mAd560_1 CB@11_mAd560_2 CB@11_mAd561_1 CB@11_mAd561_2 CB@11_mAd562_1 CB@11_mAd562_2 CB@11_mAd563_1 CB@11_mAd563_2 CB@11_mAd564_1 CB@11_mAd564_2 CB@11_mAd565_1 CB@11_mAd565_2 CB@11_mAd566_1 
+CB@11_mAd566_2 CB@11_mAd567_1 CB@11_mAd567_2 CB@11_mAd570_1 CB@11_mAd570_2 CB@11_mAd571_1 CB@11_mAd571_2 CB@11_mAd572_1 CB@11_mAd572_2 CB@11_mAd573_1 CB@11_mAd573_2 CB@11_mAd575_1 CB@11_mAd575_2 CB@11_mAd576_1 CB@11_mAd576_2 CB@11_mAd577_1 CB@11_mAd577_2 CB@11_mAd600_1 CB@11_mAd600_2 CB@11_mAd601_1 CB@11_mAd601_2 CB@11_mAd602_1 CB@11_mAd602_2 CB@11_mAd604_1 CB@11_mAd604_2 CB@11_mAd605_1 CB@11_mAd605_2 CB@11_mAd606_1 CB@11_mAd606_2 CB@11_mAd607_1 CB@11_mAd607_2 CB@11_mAd610_1 CB@11_mAd610_2 CB@11_mAd611_1 
+CB@11_mAd611_2 CB@11_mAd612_1 CB@11_mAd612_2 CB@11_mAd613_1 CB@11_mAd613_2 CB@11_mAd614_1 CB@11_mAd614_2 CB@11_mAd615_1 CB@11_mAd615_2 CB@11_mAd616_1 CB@11_mAd616_2 CB@11_mAd617_1 CB@11_mAd617_2 CB@11_mAd620_1 CB@11_mAd620_2 CB@11_mAd621_1 CB@11_mAd621_2 CB@11_mAd622_1 CB@11_mAd622_2 CB@11_mAd623_1 CB@11_mAd623_2 CB@11_mAd624_1 CB@11_mAd624_2 CB@11_mAd625_1 CB@11_mAd625_2 CB@11_mAd626_1 CB@11_mAd626_2 CB@11_mAd627_1 CB@11_mAd627_2 CB@11_mAd630_1 CB@11_mAd630_2 CB@11_mAd631_1 CB@11_mAd631_2 CB@11_mAd632_1 
+CB@11_mAd632_2 CB@11_mAd633_1 CB@11_mAd633_2 CB@11_mAd634_1 CB@11_mAd634_2 CB@11_mAd635_1 CB@11_mAd635_2 CB@11_mAd636_1 CB@11_mAd636_2 CB@11_mAd637_1 CB@11_mAd637_2 CB@11_mAd640_1 CB@11_mAd640_2 CB@11_mAd641_1 CB@11_mAd641_2 CB@11_mAd642_1 CB@11_mAd642_2 CB@11_mAd643_1 CB@11_mAd643_2 CB@11_mAd644_1 CB@11_mAd644_2 CB@11_mAd645_1 CB@11_mAd645_2 CB@11_mAd646_1 CB@11_mAd646_2 CB@11_mAd647_1 CB@11_mAd647_2 CB@11_mAd650_1 CB@11_mAd650_2 CB@11_mAd651_1 CB@11_mAd651_2 CB@11_mAd652_1 CB@11_mAd652_2 CB@11_mAd653_1 
+CB@11_mAd653_2 CB@11_mAd654_1 CB@11_mAd654_2 CB@11_mAd655_1 CB@11_mAd655_2 CB@11_mAd656_1 CB@11_mAd656_2 CB@11_mAd657_1 CB@11_mAd657_2 CB@11_mAd660_1 CB@11_mAd660_2 CB@11_mAd661_1 CB@11_mAd661_2 CB@11_mAd662_1 CB@11_mAd662_2 CB@11_mAd663_1 CB@11_mAd663_2 CB@11_mAd664_1 CB@11_mAd664_2 CB@11_mAd665_1 CB@11_mAd665_2 CB@11_mAd666_1 CB@11_mAd666_2 CB@11_mAd667_1 CB@11_mAd667_2 CB@11_mAd675_1 CB@11_mAd675_2 CB@11_mAd676_1 CB@11_mAd676_2 CB@11_mAd677_1 CB@11_mAd677_2 CB@11_mAd700_1 CB@11_mAd700_2 CB@11_mAd710_1 
+CB@11_mAd710_2 CB@11_mAd711_1 CB@11_mAd711_2 CB@11_mAd717_1 CB@11_mAd717_2 CB@11_mAd720_1 CB@11_mAd720_2 CB@11_mAd721_1 CB@11_mAd721_2 CB@11_mAd722_1 CB@11_mAd722_2 CB@11_mAd723_1 CB@11_mAd723_2 CB@11_mAd724_1 CB@11_mAd724_2 CB@11_mAd725_1 CB@11_mAd725_2 CB@11_mAd726_1 CB@11_mAd726_2 CB@11_mAd727_1 CB@11_mAd727_2 CB@11_mAd730_1 CB@11_mAd730_2 CB@11_mAd731_1 CB@11_mAd731_2 CB@11_mAd732_1 CB@11_mAd732_2 CB@11_mAd733_1 CB@11_mAd733_2 CB@11_mAd734_1 CB@11_mAd734_2 CB@11_mAd735_1 CB@11_mAd735_2 CB@11_mAd736_1 
+CB@11_mAd736_2 CB@11_mAd737_1 CB@11_mAd737_2 CB@11_mAd740_1 CB@11_mAd740_2 CB@11_mAd741_1 CB@11_mAd741_2 CB@11_mAd742_1 CB@11_mAd742_2 CB@11_mAd743_1 CB@11_mAd743_2 CB@11_mAd744_1 CB@11_mAd744_2 CB@11_mAd745_1 CB@11_mAd745_2 CB@11_mAd746_1 CB@11_mAd746_2 CB@11_mAd747_1 CB@11_mAd747_2 CB@11_mAd750_1 CB@11_mAd750_2 CB@11_mAd751_1 CB@11_mAd751_2 CB@11_mAd752_1 CB@11_mAd752_2 CB@11_mAd753_1 CB@11_mAd753_2 CB@11_mAd754_1 CB@11_mAd754_2 CB@11_mAd755_1 CB@11_mAd755_2 CB@11_mAd756_1 CB@11_mAd756_2 CB@11_mAd757_1 
+CB@11_mAd757_2 CB@11_mAd760_1 CB@11_mAd760_2 CB@11_mAd761_1 CB@11_mAd761_2 CB@11_mAd762_1 CB@11_mAd762_2 CB@11_mAd763_1 CB@11_mAd763_2 CB@11_mAd764_1 CB@11_mAd764_2 CB@11_mAd765_1 CB@11_mAd765_2 CB@11_mAd766_1 CB@11_mAd766_2 CB@11_mAd767_1 CB@11_mAd767_2 CB@11_mAd771_1 CB@11_mAd771_2 CB@11_mAd772_1 CB@11_mAd772_2 CB@11_mAd773_1 CB@11_mAd773_2 CB@11_mAd774_1 CB@11_mAd774_2 CB@11_mAd775_1 CB@11_mAd775_2 CB@11_mAd776_1 CB@11_mAd776_2 CB@11_mAd777_1 CB@11_mAd777_2 CB@11_X0 CB@11_X1 CB@11_X10 CB@11_X11 
+CB@11_X12 CB@11_X13 CB@11_X2 CB@11_X3 CB@11_X4 CB@11_X5 CB@11_X6 CB@11_X7 CB@11_X8 CB@11_X9 CB@11_Y1 CB@11_Y10 CB@11_Y11 CB@11_Y12 CB@11_Y2 CB@11_Y3 CB@11_Y4 CB@11_Y5 CB@11_Y6 CB@11_Y7 CB@11_Y8 CB@11_Y9 CB@11_Z1 CB@11_Z10 CB@11_Z11 CB@11_Z12 CB@11_Z2 CB@11_Z3 CB@11_Z4 CB@11_Z5 CB@11_Z6 CB@11_Z7 CB@11_Z8 CB@11_Z9 _5400TP094__CB
XCB@12 CB@12_K0 CB@12_K1 CB@12_K10 CB@12_K11 CB@12_K12 CB@12_K13 CB@12_K2 CB@12_K3 CB@12_K4 CB@12_K5 CB@12_K6 CB@12_K7 CB@12_K8 CB@12_K9 CB@12_mAd000_1 CB@12_mAd000_2 CB@12_mAd001_1 CB@12_mAd001_2 CB@12_mAd002_1 CB@12_mAd002_2 CB@12_mAd003_1 CB@12_mAd003_2 CB@12_mAd004_1 CB@12_mAd004_2 CB@12_mAd005_1 CB@12_mAd005_2 CB@12_mAd006_1 CB@12_mAd006_2 CB@12_mAd007_1 CB@12_mAd007_2 CB@12_mAd010_1 CB@12_mAd010_2 CB@12_mAd011_1 CB@12_mAd011_2 CB@12_mAd012_1 CB@12_mAd012_2 CB@12_mAd013_1 CB@12_mAd013_2 CB@12_mAd014_1 
+CB@12_mAd014_2 CB@12_mAd015_1 CB@12_mAd015_2 CB@12_mAd016_1 CB@12_mAd016_2 CB@12_mAd017_1 CB@12_mAd017_2 CB@12_mAd020_1 CB@12_mAd020_2 CB@12_mAd021_1 CB@12_mAd021_2 CB@12_mAd022_1 CB@12_mAd022_2 CB@12_mAd023_1 CB@12_mAd023_2 CB@12_mAd024_1 CB@12_mAd024_2 CB@12_mAd025_1 CB@12_mAd025_2 CB@12_mAd026_1 CB@12_mAd026_2 CB@12_mAd027_1 CB@12_mAd027_2 CB@12_mAd030_1 CB@12_mAd030_2 CB@12_mAd031_1 CB@12_mAd031_2 CB@12_mAd032_1 CB@12_mAd032_2 CB@12_mAd033_1 CB@12_mAd033_2 CB@12_mAd034_1 CB@12_mAd034_2 CB@12_mAd035_1 
+CB@12_mAd035_2 CB@12_mAd036_1 CB@12_mAd036_2 CB@12_mAd037_1 CB@12_mAd037_2 CB@12_mAd040_1 CB@12_mAd040_2 CB@12_mAd041_1 CB@12_mAd041_2 CB@12_mAd042_1 CB@12_mAd042_2 CB@12_mAd043_1 CB@12_mAd043_2 CB@12_mAd044_1 CB@12_mAd044_2 CB@12_mAd045_1 CB@12_mAd045_2 CB@12_mAd046_1 CB@12_mAd046_2 CB@12_mAd047_1 CB@12_mAd047_2 CB@12_mAd050_1 CB@12_mAd050_2 CB@12_mAd051_1 CB@12_mAd051_2 CB@12_mAd052_1 CB@12_mAd052_2 CB@12_mAd053_1 CB@12_mAd053_2 CB@12_mAd054_1 CB@12_mAd054_2 CB@12_mAd055_1 CB@12_mAd055_2 CB@12_mAd056_1 
+CB@12_mAd056_2 CB@12_mAd057_1 CB@12_mAd057_2 CB@12_mAd060_1 CB@12_mAd060_2 CB@12_mAd066_1 CB@12_mAd066_2 CB@12_mAd067_1 CB@12_mAd067_2 CB@12_mAd100_1 CB@12_mAd100_2 CB@12_mAd101_1 CB@12_mAd101_2 CB@12_mAd102_1 CB@12_mAd102_2 CB@12_mAd110_1 CB@12_mAd110_2 CB@12_mAd111_1 CB@12_mAd111_2 CB@12_mAd112_1 CB@12_mAd112_2 CB@12_mAd113_1 CB@12_mAd113_2 CB@12_mAd114_1 CB@12_mAd114_2 CB@12_mAd115_1 CB@12_mAd115_2 CB@12_mAd116_1 CB@12_mAd116_2 CB@12_mAd117_1 CB@12_mAd117_2 CB@12_mAd120_1 CB@12_mAd120_2 CB@12_mAd121_1 
+CB@12_mAd121_2 CB@12_mAd122_1 CB@12_mAd122_2 CB@12_mAd123_1 CB@12_mAd123_2 CB@12_mAd124_1 CB@12_mAd124_2 CB@12_mAd125_1 CB@12_mAd125_2 CB@12_mAd126_1 CB@12_mAd126_2 CB@12_mAd127_1 CB@12_mAd127_2 CB@12_mAd130_1 CB@12_mAd130_2 CB@12_mAd131_1 CB@12_mAd131_2 CB@12_mAd132_1 CB@12_mAd132_2 CB@12_mAd133_1 CB@12_mAd133_2 CB@12_mAd134_1 CB@12_mAd134_2 CB@12_mAd135_1 CB@12_mAd135_2 CB@12_mAd136_1 CB@12_mAd136_2 CB@12_mAd137_1 CB@12_mAd137_2 CB@12_mAd140_1 CB@12_mAd140_2 CB@12_mAd141_1 CB@12_mAd141_2 CB@12_mAd142_1 
+CB@12_mAd142_2 CB@12_mAd143_1 CB@12_mAd143_2 CB@12_mAd144_1 CB@12_mAd144_2 CB@12_mAd145_1 CB@12_mAd145_2 CB@12_mAd146_1 CB@12_mAd146_2 CB@12_mAd147_1 CB@12_mAd147_2 CB@12_mAd150_1 CB@12_mAd150_2 CB@12_mAd151_1 CB@12_mAd151_2 CB@12_mAd152_1 CB@12_mAd152_2 CB@12_mAd153_1 CB@12_mAd153_2 CB@12_mAd154_1 CB@12_mAd154_2 CB@12_mAd155_1 CB@12_mAd155_2 CB@12_mAd156_1 CB@12_mAd156_2 CB@12_mAd157_1 CB@12_mAd157_2 CB@12_mAd160_1 CB@12_mAd160_2 CB@12_mAd161_1 CB@12_mAd161_2 CB@12_mAd162_1 CB@12_mAd162_2 CB@12_mAd163_1 
+CB@12_mAd163_2 CB@12_mAd164_1 CB@12_mAd164_2 CB@12_mAd165_1 CB@12_mAd165_2 CB@12_mAd166_1 CB@12_mAd166_2 CB@12_mAd167_1 CB@12_mAd167_2 CB@12_mAd170_1 CB@12_mAd170_2 CB@12_mAd171_1 CB@12_mAd171_2 CB@12_mAd172_1 CB@12_mAd172_2 CB@12_mAd173_1 CB@12_mAd173_2 CB@12_mAd175_1 CB@12_mAd175_2 CB@12_mAd176_1 CB@12_mAd176_2 CB@12_mAd177_1 CB@12_mAd177_2 CB@12_mAd200_1 CB@12_mAd200_2 CB@12_mAd201_1 CB@12_mAd201_2 CB@12_mAd202_1 CB@12_mAd202_2 CB@12_mAd204_1 CB@12_mAd204_2 CB@12_mAd205_1 CB@12_mAd205_2 CB@12_mAd206_1 
+CB@12_mAd206_2 CB@12_mAd207_1 CB@12_mAd207_2 CB@12_mAd210_1 CB@12_mAd210_2 CB@12_mAd211_1 CB@12_mAd211_2 CB@12_mAd212_1 CB@12_mAd212_2 CB@12_mAd213_1 CB@12_mAd213_2 CB@12_mAd214_1 CB@12_mAd214_2 CB@12_mAd215_1 CB@12_mAd215_2 CB@12_mAd216_1 CB@12_mAd216_2 CB@12_mAd217_1 CB@12_mAd217_2 CB@12_mAd220_1 CB@12_mAd220_2 CB@12_mAd221_1 CB@12_mAd221_2 CB@12_mAd222_1 CB@12_mAd222_2 CB@12_mAd223_1 CB@12_mAd223_2 CB@12_mAd224_1 CB@12_mAd224_2 CB@12_mAd225_1 CB@12_mAd225_2 CB@12_mAd226_1 CB@12_mAd226_2 CB@12_mAd227_1 
+CB@12_mAd227_2 CB@12_mAd230_1 CB@12_mAd230_2 CB@12_mAd231_1 CB@12_mAd231_2 CB@12_mAd232_1 CB@12_mAd232_2 CB@12_mAd233_1 CB@12_mAd233_2 CB@12_mAd234_1 CB@12_mAd234_2 CB@12_mAd235_1 CB@12_mAd235_2 CB@12_mAd236_1 CB@12_mAd236_2 CB@12_mAd237_1 CB@12_mAd237_2 CB@12_mAd240_1 CB@12_mAd240_2 CB@12_mAd241_1 CB@12_mAd241_2 CB@12_mAd242_1 CB@12_mAd242_2 CB@12_mAd243_1 CB@12_mAd243_2 CB@12_mAd244_1 CB@12_mAd244_2 CB@12_mAd245_1 CB@12_mAd245_2 CB@12_mAd246_1 CB@12_mAd246_2 CB@12_mAd247_1 CB@12_mAd247_2 CB@12_mAd250_1 
+CB@12_mAd250_2 CB@12_mAd251_1 CB@12_mAd251_2 CB@12_mAd252_1 CB@12_mAd252_2 CB@12_mAd253_1 CB@12_mAd253_2 CB@12_mAd254_1 CB@12_mAd254_2 CB@12_mAd255_1 CB@12_mAd255_2 CB@12_mAd256_1 CB@12_mAd256_2 CB@12_mAd257_1 CB@12_mAd257_2 CB@12_mAd260_1 CB@12_mAd260_2 CB@12_mAd261_1 CB@12_mAd261_2 CB@12_mAd262_1 CB@12_mAd262_2 CB@12_mAd263_1 CB@12_mAd263_2 CB@12_mAd264_1 CB@12_mAd264_2 CB@12_mAd265_1 CB@12_mAd265_2 CB@12_mAd266_1 CB@12_mAd266_2 CB@12_mAd267_1 CB@12_mAd267_2 CB@12_mAd275_1 CB@12_mAd275_2 CB@12_mAd276_1 
+CB@12_mAd276_2 CB@12_mAd277_1 CB@12_mAd277_2 CB@12_mAd300_1 CB@12_mAd300_2 CB@12_mAd310_1 CB@12_mAd310_2 CB@12_mAd311_1 CB@12_mAd311_2 CB@12_mAd317_1 CB@12_mAd317_2 CB@12_mAd320_1 CB@12_mAd320_2 CB@12_mAd321_1 CB@12_mAd321_2 CB@12_mAd322_1 CB@12_mAd322_2 CB@12_mAd323_1 CB@12_mAd323_2 CB@12_mAd324_1 CB@12_mAd324_2 CB@12_mAd325_1 CB@12_mAd325_2 CB@12_mAd326_1 CB@12_mAd326_2 CB@12_mAd327_1 CB@12_mAd327_2 CB@12_mAd330_1 CB@12_mAd330_2 CB@12_mAd331_1 CB@12_mAd331_2 CB@12_mAd332_1 CB@12_mAd332_2 CB@12_mAd333_1 
+CB@12_mAd333_2 CB@12_mAd334_1 CB@12_mAd334_2 CB@12_mAd335_1 CB@12_mAd335_2 CB@12_mAd336_1 CB@12_mAd336_2 CB@12_mAd337_1 CB@12_mAd337_2 CB@12_mAd340_1 CB@12_mAd340_2 CB@12_mAd341_1 CB@12_mAd341_2 CB@12_mAd342_1 CB@12_mAd342_2 CB@12_mAd343_1 CB@12_mAd343_2 CB@12_mAd344_1 CB@12_mAd344_2 CB@12_mAd345_1 CB@12_mAd345_2 CB@12_mAd346_1 CB@12_mAd346_2 CB@12_mAd347_1 CB@12_mAd347_2 CB@12_mAd350_1 CB@12_mAd350_2 CB@12_mAd351_1 CB@12_mAd351_2 CB@12_mAd352_1 CB@12_mAd352_2 CB@12_mAd353_1 CB@12_mAd353_2 CB@12_mAd354_1 
+CB@12_mAd354_2 CB@12_mAd355_1 CB@12_mAd355_2 CB@12_mAd356_1 CB@12_mAd356_2 CB@12_mAd357_1 CB@12_mAd357_2 CB@12_mAd360_1 CB@12_mAd360_2 CB@12_mAd361_1 CB@12_mAd361_2 CB@12_mAd362_1 CB@12_mAd362_2 CB@12_mAd363_1 CB@12_mAd363_2 CB@12_mAd364_1 CB@12_mAd364_2 CB@12_mAd365_1 CB@12_mAd365_2 CB@12_mAd366_1 CB@12_mAd366_2 CB@12_mAd367_1 CB@12_mAd367_2 CB@12_mAd371_1 CB@12_mAd371_2 CB@12_mAd372_1 CB@12_mAd372_2 CB@12_mAd373_1 CB@12_mAd373_2 CB@12_mAd374_1 CB@12_mAd374_2 CB@12_mAd375_1 CB@12_mAd375_2 CB@12_mAd376_1 
+CB@12_mAd376_2 CB@12_mAd377_1 CB@12_mAd377_2 CB@12_mAd400_1 CB@12_mAd400_2 CB@12_mAd401_1 CB@12_mAd401_2 CB@12_mAd402_1 CB@12_mAd402_2 CB@12_mAd403_1 CB@12_mAd403_2 CB@12_mAd404_1 CB@12_mAd404_2 CB@12_mAd405_1 CB@12_mAd405_2 CB@12_mAd406_1 CB@12_mAd406_2 CB@12_mAd407_1 CB@12_mAd407_2 CB@12_mAd410_1 CB@12_mAd410_2 CB@12_mAd411_1 CB@12_mAd411_2 CB@12_mAd412_1 CB@12_mAd412_2 CB@12_mAd413_1 CB@12_mAd413_2 CB@12_mAd414_1 CB@12_mAd414_2 CB@12_mAd415_1 CB@12_mAd415_2 CB@12_mAd416_1 CB@12_mAd416_2 CB@12_mAd417_1 
+CB@12_mAd417_2 CB@12_mAd420_1 CB@12_mAd420_2 CB@12_mAd421_1 CB@12_mAd421_2 CB@12_mAd422_1 CB@12_mAd422_2 CB@12_mAd423_1 CB@12_mAd423_2 CB@12_mAd424_1 CB@12_mAd424_2 CB@12_mAd425_1 CB@12_mAd425_2 CB@12_mAd426_1 CB@12_mAd426_2 CB@12_mAd427_1 CB@12_mAd427_2 CB@12_mAd430_1 CB@12_mAd430_2 CB@12_mAd431_1 CB@12_mAd431_2 CB@12_mAd432_1 CB@12_mAd432_2 CB@12_mAd433_1 CB@12_mAd433_2 CB@12_mAd434_1 CB@12_mAd434_2 CB@12_mAd435_1 CB@12_mAd435_2 CB@12_mAd436_1 CB@12_mAd436_2 CB@12_mAd437_1 CB@12_mAd437_2 CB@12_mAd440_1 
+CB@12_mAd440_2 CB@12_mAd441_1 CB@12_mAd441_2 CB@12_mAd442_1 CB@12_mAd442_2 CB@12_mAd443_1 CB@12_mAd443_2 CB@12_mAd444_1 CB@12_mAd444_2 CB@12_mAd445_1 CB@12_mAd445_2 CB@12_mAd446_1 CB@12_mAd446_2 CB@12_mAd447_1 CB@12_mAd447_2 CB@12_mAd450_1 CB@12_mAd450_2 CB@12_mAd451_1 CB@12_mAd451_2 CB@12_mAd452_1 CB@12_mAd452_2 CB@12_mAd453_1 CB@12_mAd453_2 CB@12_mAd454_1 CB@12_mAd454_2 CB@12_mAd455_1 CB@12_mAd455_2 CB@12_mAd456_1 CB@12_mAd456_2 CB@12_mAd457_1 CB@12_mAd457_2 CB@12_mAd460_1 CB@12_mAd460_2 CB@12_mAd466_1 
+CB@12_mAd466_2 CB@12_mAd467_1 CB@12_mAd467_2 CB@12_mAd500_1 CB@12_mAd500_2 CB@12_mAd501_1 CB@12_mAd501_2 CB@12_mAd502_1 CB@12_mAd502_2 CB@12_mAd508_1 CB@12_mAd508_2 CB@12_mAd509_1 CB@12_mAd509_2 CB@12_mAd512_1 CB@12_mAd512_2 CB@12_mAd513_1 CB@12_mAd513_2 CB@12_mAd514_1 CB@12_mAd514_2 CB@12_mAd515_1 CB@12_mAd515_2 CB@12_mAd516_1 CB@12_mAd516_2 CB@12_mAd517_1 CB@12_mAd517_2 CB@12_mAd520_1 CB@12_mAd520_2 CB@12_mAd521_1 CB@12_mAd521_2 CB@12_mAd522_1 CB@12_mAd522_2 CB@12_mAd523_1 CB@12_mAd523_2 CB@12_mAd524_1 
+CB@12_mAd524_2 CB@12_mAd525_1 CB@12_mAd525_2 CB@12_mAd526_1 CB@12_mAd526_2 CB@12_mAd527_1 CB@12_mAd527_2 CB@12_mAd530_1 CB@12_mAd530_2 CB@12_mAd531_1 CB@12_mAd531_2 CB@12_mAd532_1 CB@12_mAd532_2 CB@12_mAd533_1 CB@12_mAd533_2 CB@12_mAd534_1 CB@12_mAd534_2 CB@12_mAd535_1 CB@12_mAd535_2 CB@12_mAd536_1 CB@12_mAd536_2 CB@12_mAd537_1 CB@12_mAd537_2 CB@12_mAd540_1 CB@12_mAd540_2 CB@12_mAd541_1 CB@12_mAd541_2 CB@12_mAd542_1 CB@12_mAd542_2 CB@12_mAd543_1 CB@12_mAd543_2 CB@12_mAd544_1 CB@12_mAd544_2 CB@12_mAd545_1 
+CB@12_mAd545_2 CB@12_mAd546_1 CB@12_mAd546_2 CB@12_mAd547_1 CB@12_mAd547_2 CB@12_mAd550_1 CB@12_mAd550_2 CB@12_mAd551_1 CB@12_mAd551_2 CB@12_mAd552_1 CB@12_mAd552_2 CB@12_mAd553_1 CB@12_mAd553_2 CB@12_mAd554_1 CB@12_mAd554_2 CB@12_mAd555_1 CB@12_mAd555_2 CB@12_mAd556_1 CB@12_mAd556_2 CB@12_mAd557_1 CB@12_mAd557_2 CB@12_mAd560_1 CB@12_mAd560_2 CB@12_mAd561_1 CB@12_mAd561_2 CB@12_mAd562_1 CB@12_mAd562_2 CB@12_mAd563_1 CB@12_mAd563_2 CB@12_mAd564_1 CB@12_mAd564_2 CB@12_mAd565_1 CB@12_mAd565_2 CB@12_mAd566_1 
+CB@12_mAd566_2 CB@12_mAd567_1 CB@12_mAd567_2 CB@12_mAd570_1 CB@12_mAd570_2 CB@12_mAd571_1 CB@12_mAd571_2 CB@12_mAd572_1 CB@12_mAd572_2 CB@12_mAd573_1 CB@12_mAd573_2 CB@12_mAd575_1 CB@12_mAd575_2 CB@12_mAd576_1 CB@12_mAd576_2 CB@12_mAd577_1 CB@12_mAd577_2 CB@12_mAd600_1 CB@12_mAd600_2 CB@12_mAd601_1 CB@12_mAd601_2 CB@12_mAd602_1 CB@12_mAd602_2 CB@12_mAd604_1 CB@12_mAd604_2 CB@12_mAd605_1 CB@12_mAd605_2 CB@12_mAd606_1 CB@12_mAd606_2 CB@12_mAd607_1 CB@12_mAd607_2 CB@12_mAd610_1 CB@12_mAd610_2 CB@12_mAd611_1 
+CB@12_mAd611_2 CB@12_mAd612_1 CB@12_mAd612_2 CB@12_mAd613_1 CB@12_mAd613_2 CB@12_mAd614_1 CB@12_mAd614_2 CB@12_mAd615_1 CB@12_mAd615_2 CB@12_mAd616_1 CB@12_mAd616_2 CB@12_mAd617_1 CB@12_mAd617_2 CB@12_mAd620_1 CB@12_mAd620_2 CB@12_mAd621_1 CB@12_mAd621_2 CB@12_mAd622_1 CB@12_mAd622_2 CB@12_mAd623_1 CB@12_mAd623_2 CB@12_mAd624_1 CB@12_mAd624_2 CB@12_mAd625_1 CB@12_mAd625_2 CB@12_mAd626_1 CB@12_mAd626_2 CB@12_mAd627_1 CB@12_mAd627_2 CB@12_mAd630_1 CB@12_mAd630_2 CB@12_mAd631_1 CB@12_mAd631_2 CB@12_mAd632_1 
+CB@12_mAd632_2 CB@12_mAd633_1 CB@12_mAd633_2 CB@12_mAd634_1 CB@12_mAd634_2 CB@12_mAd635_1 CB@12_mAd635_2 CB@12_mAd636_1 CB@12_mAd636_2 CB@12_mAd637_1 CB@12_mAd637_2 CB@12_mAd640_1 CB@12_mAd640_2 CB@12_mAd641_1 CB@12_mAd641_2 CB@12_mAd642_1 CB@12_mAd642_2 CB@12_mAd643_1 CB@12_mAd643_2 CB@12_mAd644_1 CB@12_mAd644_2 CB@12_mAd645_1 CB@12_mAd645_2 CB@12_mAd646_1 CB@12_mAd646_2 CB@12_mAd647_1 CB@12_mAd647_2 CB@12_mAd650_1 CB@12_mAd650_2 CB@12_mAd651_1 CB@12_mAd651_2 CB@12_mAd652_1 CB@12_mAd652_2 CB@12_mAd653_1 
+CB@12_mAd653_2 CB@12_mAd654_1 CB@12_mAd654_2 CB@12_mAd655_1 CB@12_mAd655_2 CB@12_mAd656_1 CB@12_mAd656_2 CB@12_mAd657_1 CB@12_mAd657_2 CB@12_mAd660_1 CB@12_mAd660_2 CB@12_mAd661_1 CB@12_mAd661_2 CB@12_mAd662_1 CB@12_mAd662_2 CB@12_mAd663_1 CB@12_mAd663_2 CB@12_mAd664_1 CB@12_mAd664_2 CB@12_mAd665_1 CB@12_mAd665_2 CB@12_mAd666_1 CB@12_mAd666_2 CB@12_mAd667_1 CB@12_mAd667_2 CB@12_mAd675_1 CB@12_mAd675_2 CB@12_mAd676_1 CB@12_mAd676_2 CB@12_mAd677_1 CB@12_mAd677_2 CB@12_mAd700_1 CB@12_mAd700_2 CB@12_mAd710_1 
+CB@12_mAd710_2 CB@12_mAd711_1 CB@12_mAd711_2 CB@12_mAd717_1 CB@12_mAd717_2 CB@12_mAd720_1 CB@12_mAd720_2 CB@12_mAd721_1 CB@12_mAd721_2 CB@12_mAd722_1 CB@12_mAd722_2 CB@12_mAd723_1 CB@12_mAd723_2 CB@12_mAd724_1 CB@12_mAd724_2 CB@12_mAd725_1 CB@12_mAd725_2 CB@12_mAd726_1 CB@12_mAd726_2 CB@12_mAd727_1 CB@12_mAd727_2 CB@12_mAd730_1 CB@12_mAd730_2 CB@12_mAd731_1 CB@12_mAd731_2 CB@12_mAd732_1 CB@12_mAd732_2 CB@12_mAd733_1 CB@12_mAd733_2 CB@12_mAd734_1 CB@12_mAd734_2 CB@12_mAd735_1 CB@12_mAd735_2 CB@12_mAd736_1 
+CB@12_mAd736_2 CB@12_mAd737_1 CB@12_mAd737_2 CB@12_mAd740_1 CB@12_mAd740_2 CB@12_mAd741_1 CB@12_mAd741_2 CB@12_mAd742_1 CB@12_mAd742_2 CB@12_mAd743_1 CB@12_mAd743_2 CB@12_mAd744_1 CB@12_mAd744_2 CB@12_mAd745_1 CB@12_mAd745_2 CB@12_mAd746_1 CB@12_mAd746_2 CB@12_mAd747_1 CB@12_mAd747_2 CB@12_mAd750_1 CB@12_mAd750_2 CB@12_mAd751_1 CB@12_mAd751_2 CB@12_mAd752_1 CB@12_mAd752_2 CB@12_mAd753_1 CB@12_mAd753_2 CB@12_mAd754_1 CB@12_mAd754_2 CB@12_mAd755_1 CB@12_mAd755_2 CB@12_mAd756_1 CB@12_mAd756_2 CB@12_mAd757_1 
+CB@12_mAd757_2 CB@12_mAd760_1 CB@12_mAd760_2 CB@12_mAd761_1 CB@12_mAd761_2 CB@12_mAd762_1 CB@12_mAd762_2 CB@12_mAd763_1 CB@12_mAd763_2 CB@12_mAd764_1 CB@12_mAd764_2 CB@12_mAd765_1 CB@12_mAd765_2 CB@12_mAd766_1 CB@12_mAd766_2 CB@12_mAd767_1 CB@12_mAd767_2 CB@12_mAd771_1 CB@12_mAd771_2 CB@12_mAd772_1 CB@12_mAd772_2 CB@12_mAd773_1 CB@12_mAd773_2 CB@12_mAd774_1 CB@12_mAd774_2 CB@12_mAd775_1 CB@12_mAd775_2 CB@12_mAd776_1 CB@12_mAd776_2 CB@12_mAd777_1 CB@12_mAd777_2 CB@12_X0 CB@12_X1 CB@12_X10 CB@12_X11 
+CB@12_X12 CB@12_X13 CB@12_X2 CB@12_X3 CB@12_X4 CB@12_X5 CB@12_X6 CB@12_X7 CB@12_X8 CB@12_X9 CB@12_Y1 CB@12_Y10 CB@12_Y11 CB@12_Y12 CB@12_Y2 CB@12_Y3 CB@12_Y4 CB@12_Y5 CB@12_Y6 CB@12_Y7 CB@12_Y8 CB@12_Y9 CB@12_Z1 CB@12_Z10 CB@12_Z11 CB@12_Z12 CB@12_Z2 CB@12_Z3 CB@12_Z4 CB@12_Z5 CB@12_Z6 CB@12_Z7 CB@12_Z8 CB@12_Z9 _5400TP094__CB
XCB@13 CB@13_K0 CB@13_K1 CB@13_K10 CB@13_K11 CB@13_K12 CB@13_K13 CB@13_K2 CB@13_K3 CB@13_K4 CB@13_K5 CB@13_K6 CB@13_K7 CB@13_K8 CB@13_K9 CB@13_mAd000_1 CB@13_mAd000_2 CB@13_mAd001_1 CB@13_mAd001_2 CB@13_mAd002_1 CB@13_mAd002_2 CB@13_mAd003_1 CB@13_mAd003_2 CB@13_mAd004_1 CB@13_mAd004_2 CB@13_mAd005_1 CB@13_mAd005_2 CB@13_mAd006_1 CB@13_mAd006_2 CB@13_mAd007_1 CB@13_mAd007_2 CB@13_mAd010_1 CB@13_mAd010_2 CB@13_mAd011_1 CB@13_mAd011_2 CB@13_mAd012_1 CB@13_mAd012_2 CB@13_mAd013_1 CB@13_mAd013_2 CB@13_mAd014_1 
+CB@13_mAd014_2 CB@13_mAd015_1 CB@13_mAd015_2 CB@13_mAd016_1 CB@13_mAd016_2 CB@13_mAd017_1 CB@13_mAd017_2 CB@13_mAd020_1 CB@13_mAd020_2 CB@13_mAd021_1 CB@13_mAd021_2 CB@13_mAd022_1 CB@13_mAd022_2 CB@13_mAd023_1 CB@13_mAd023_2 CB@13_mAd024_1 CB@13_mAd024_2 CB@13_mAd025_1 CB@13_mAd025_2 CB@13_mAd026_1 CB@13_mAd026_2 CB@13_mAd027_1 CB@13_mAd027_2 CB@13_mAd030_1 CB@13_mAd030_2 CB@13_mAd031_1 CB@13_mAd031_2 CB@13_mAd032_1 CB@13_mAd032_2 CB@13_mAd033_1 CB@13_mAd033_2 CB@13_mAd034_1 CB@13_mAd034_2 CB@13_mAd035_1 
+CB@13_mAd035_2 CB@13_mAd036_1 CB@13_mAd036_2 CB@13_mAd037_1 CB@13_mAd037_2 CB@13_mAd040_1 CB@13_mAd040_2 CB@13_mAd041_1 CB@13_mAd041_2 CB@13_mAd042_1 CB@13_mAd042_2 CB@13_mAd043_1 CB@13_mAd043_2 CB@13_mAd044_1 CB@13_mAd044_2 CB@13_mAd045_1 CB@13_mAd045_2 CB@13_mAd046_1 CB@13_mAd046_2 CB@13_mAd047_1 CB@13_mAd047_2 CB@13_mAd050_1 CB@13_mAd050_2 CB@13_mAd051_1 CB@13_mAd051_2 CB@13_mAd052_1 CB@13_mAd052_2 CB@13_mAd053_1 CB@13_mAd053_2 CB@13_mAd054_1 CB@13_mAd054_2 CB@13_mAd055_1 CB@13_mAd055_2 CB@13_mAd056_1 
+CB@13_mAd056_2 CB@13_mAd057_1 CB@13_mAd057_2 CB@13_mAd060_1 CB@13_mAd060_2 CB@13_mAd066_1 CB@13_mAd066_2 CB@13_mAd067_1 CB@13_mAd067_2 CB@13_mAd100_1 CB@13_mAd100_2 CB@13_mAd101_1 CB@13_mAd101_2 CB@13_mAd102_1 CB@13_mAd102_2 CB@13_mAd110_1 CB@13_mAd110_2 CB@13_mAd111_1 CB@13_mAd111_2 CB@13_mAd112_1 CB@13_mAd112_2 CB@13_mAd113_1 CB@13_mAd113_2 CB@13_mAd114_1 CB@13_mAd114_2 CB@13_mAd115_1 CB@13_mAd115_2 CB@13_mAd116_1 CB@13_mAd116_2 CB@13_mAd117_1 CB@13_mAd117_2 CB@13_mAd120_1 CB@13_mAd120_2 CB@13_mAd121_1 
+CB@13_mAd121_2 CB@13_mAd122_1 CB@13_mAd122_2 CB@13_mAd123_1 CB@13_mAd123_2 CB@13_mAd124_1 CB@13_mAd124_2 CB@13_mAd125_1 CB@13_mAd125_2 CB@13_mAd126_1 CB@13_mAd126_2 CB@13_mAd127_1 CB@13_mAd127_2 CB@13_mAd130_1 CB@13_mAd130_2 CB@13_mAd131_1 CB@13_mAd131_2 CB@13_mAd132_1 CB@13_mAd132_2 CB@13_mAd133_1 CB@13_mAd133_2 CB@13_mAd134_1 CB@13_mAd134_2 CB@13_mAd135_1 CB@13_mAd135_2 CB@13_mAd136_1 CB@13_mAd136_2 CB@13_mAd137_1 CB@13_mAd137_2 CB@13_mAd140_1 CB@13_mAd140_2 CB@13_mAd141_1 CB@13_mAd141_2 CB@13_mAd142_1 
+CB@13_mAd142_2 CB@13_mAd143_1 CB@13_mAd143_2 CB@13_mAd144_1 CB@13_mAd144_2 CB@13_mAd145_1 CB@13_mAd145_2 CB@13_mAd146_1 CB@13_mAd146_2 CB@13_mAd147_1 CB@13_mAd147_2 CB@13_mAd150_1 CB@13_mAd150_2 CB@13_mAd151_1 CB@13_mAd151_2 CB@13_mAd152_1 CB@13_mAd152_2 CB@13_mAd153_1 CB@13_mAd153_2 CB@13_mAd154_1 CB@13_mAd154_2 CB@13_mAd155_1 CB@13_mAd155_2 CB@13_mAd156_1 CB@13_mAd156_2 CB@13_mAd157_1 CB@13_mAd157_2 CB@13_mAd160_1 CB@13_mAd160_2 CB@13_mAd161_1 CB@13_mAd161_2 CB@13_mAd162_1 CB@13_mAd162_2 CB@13_mAd163_1 
+CB@13_mAd163_2 CB@13_mAd164_1 CB@13_mAd164_2 CB@13_mAd165_1 CB@13_mAd165_2 CB@13_mAd166_1 CB@13_mAd166_2 CB@13_mAd167_1 CB@13_mAd167_2 CB@13_mAd170_1 CB@13_mAd170_2 CB@13_mAd171_1 CB@13_mAd171_2 CB@13_mAd172_1 CB@13_mAd172_2 CB@13_mAd173_1 CB@13_mAd173_2 CB@13_mAd175_1 CB@13_mAd175_2 CB@13_mAd176_1 CB@13_mAd176_2 CB@13_mAd177_1 CB@13_mAd177_2 CB@13_mAd200_1 CB@13_mAd200_2 CB@13_mAd201_1 CB@13_mAd201_2 CB@13_mAd202_1 CB@13_mAd202_2 CB@13_mAd204_1 CB@13_mAd204_2 CB@13_mAd205_1 CB@13_mAd205_2 CB@13_mAd206_1 
+CB@13_mAd206_2 CB@13_mAd207_1 CB@13_mAd207_2 CB@13_mAd210_1 CB@13_mAd210_2 CB@13_mAd211_1 CB@13_mAd211_2 CB@13_mAd212_1 CB@13_mAd212_2 CB@13_mAd213_1 CB@13_mAd213_2 CB@13_mAd214_1 CB@13_mAd214_2 CB@13_mAd215_1 CB@13_mAd215_2 CB@13_mAd216_1 CB@13_mAd216_2 CB@13_mAd217_1 CB@13_mAd217_2 CB@13_mAd220_1 CB@13_mAd220_2 CB@13_mAd221_1 CB@13_mAd221_2 CB@13_mAd222_1 CB@13_mAd222_2 CB@13_mAd223_1 CB@13_mAd223_2 CB@13_mAd224_1 CB@13_mAd224_2 CB@13_mAd225_1 CB@13_mAd225_2 CB@13_mAd226_1 CB@13_mAd226_2 CB@13_mAd227_1 
+CB@13_mAd227_2 CB@13_mAd230_1 CB@13_mAd230_2 CB@13_mAd231_1 CB@13_mAd231_2 CB@13_mAd232_1 CB@13_mAd232_2 CB@13_mAd233_1 CB@13_mAd233_2 CB@13_mAd234_1 CB@13_mAd234_2 CB@13_mAd235_1 CB@13_mAd235_2 CB@13_mAd236_1 CB@13_mAd236_2 CB@13_mAd237_1 CB@13_mAd237_2 CB@13_mAd240_1 CB@13_mAd240_2 CB@13_mAd241_1 CB@13_mAd241_2 CB@13_mAd242_1 CB@13_mAd242_2 CB@13_mAd243_1 CB@13_mAd243_2 CB@13_mAd244_1 CB@13_mAd244_2 CB@13_mAd245_1 CB@13_mAd245_2 CB@13_mAd246_1 CB@13_mAd246_2 CB@13_mAd247_1 CB@13_mAd247_2 CB@13_mAd250_1 
+CB@13_mAd250_2 CB@13_mAd251_1 CB@13_mAd251_2 CB@13_mAd252_1 CB@13_mAd252_2 CB@13_mAd253_1 CB@13_mAd253_2 CB@13_mAd254_1 CB@13_mAd254_2 CB@13_mAd255_1 CB@13_mAd255_2 CB@13_mAd256_1 CB@13_mAd256_2 CB@13_mAd257_1 CB@13_mAd257_2 CB@13_mAd260_1 CB@13_mAd260_2 CB@13_mAd261_1 CB@13_mAd261_2 CB@13_mAd262_1 CB@13_mAd262_2 CB@13_mAd263_1 CB@13_mAd263_2 CB@13_mAd264_1 CB@13_mAd264_2 CB@13_mAd265_1 CB@13_mAd265_2 CB@13_mAd266_1 CB@13_mAd266_2 CB@13_mAd267_1 CB@13_mAd267_2 CB@13_mAd275_1 CB@13_mAd275_2 CB@13_mAd276_1 
+CB@13_mAd276_2 CB@13_mAd277_1 CB@13_mAd277_2 CB@13_mAd300_1 CB@13_mAd300_2 CB@13_mAd310_1 CB@13_mAd310_2 CB@13_mAd311_1 CB@13_mAd311_2 CB@13_mAd317_1 CB@13_mAd317_2 CB@13_mAd320_1 CB@13_mAd320_2 CB@13_mAd321_1 CB@13_mAd321_2 CB@13_mAd322_1 CB@13_mAd322_2 CB@13_mAd323_1 CB@13_mAd323_2 CB@13_mAd324_1 CB@13_mAd324_2 CB@13_mAd325_1 CB@13_mAd325_2 CB@13_mAd326_1 CB@13_mAd326_2 CB@13_mAd327_1 CB@13_mAd327_2 CB@13_mAd330_1 CB@13_mAd330_2 CB@13_mAd331_1 CB@13_mAd331_2 CB@13_mAd332_1 CB@13_mAd332_2 CB@13_mAd333_1 
+CB@13_mAd333_2 CB@13_mAd334_1 CB@13_mAd334_2 CB@13_mAd335_1 CB@13_mAd335_2 CB@13_mAd336_1 CB@13_mAd336_2 CB@13_mAd337_1 CB@13_mAd337_2 CB@13_mAd340_1 CB@13_mAd340_2 CB@13_mAd341_1 CB@13_mAd341_2 CB@13_mAd342_1 CB@13_mAd342_2 CB@13_mAd343_1 CB@13_mAd343_2 CB@13_mAd344_1 CB@13_mAd344_2 CB@13_mAd345_1 CB@13_mAd345_2 CB@13_mAd346_1 CB@13_mAd346_2 CB@13_mAd347_1 CB@13_mAd347_2 CB@13_mAd350_1 CB@13_mAd350_2 CB@13_mAd351_1 CB@13_mAd351_2 CB@13_mAd352_1 CB@13_mAd352_2 CB@13_mAd353_1 CB@13_mAd353_2 CB@13_mAd354_1 
+CB@13_mAd354_2 CB@13_mAd355_1 CB@13_mAd355_2 CB@13_mAd356_1 CB@13_mAd356_2 CB@13_mAd357_1 CB@13_mAd357_2 CB@13_mAd360_1 CB@13_mAd360_2 CB@13_mAd361_1 CB@13_mAd361_2 CB@13_mAd362_1 CB@13_mAd362_2 CB@13_mAd363_1 CB@13_mAd363_2 CB@13_mAd364_1 CB@13_mAd364_2 CB@13_mAd365_1 CB@13_mAd365_2 CB@13_mAd366_1 CB@13_mAd366_2 CB@13_mAd367_1 CB@13_mAd367_2 CB@13_mAd371_1 CB@13_mAd371_2 CB@13_mAd372_1 CB@13_mAd372_2 CB@13_mAd373_1 CB@13_mAd373_2 CB@13_mAd374_1 CB@13_mAd374_2 CB@13_mAd375_1 CB@13_mAd375_2 CB@13_mAd376_1 
+CB@13_mAd376_2 CB@13_mAd377_1 CB@13_mAd377_2 CB@13_mAd400_1 CB@13_mAd400_2 CB@13_mAd401_1 CB@13_mAd401_2 CB@13_mAd402_1 CB@13_mAd402_2 CB@13_mAd403_1 CB@13_mAd403_2 CB@13_mAd404_1 CB@13_mAd404_2 CB@13_mAd405_1 CB@13_mAd405_2 CB@13_mAd406_1 CB@13_mAd406_2 CB@13_mAd407_1 CB@13_mAd407_2 CB@13_mAd410_1 CB@13_mAd410_2 CB@13_mAd411_1 CB@13_mAd411_2 CB@13_mAd412_1 CB@13_mAd412_2 CB@13_mAd413_1 CB@13_mAd413_2 CB@13_mAd414_1 CB@13_mAd414_2 CB@13_mAd415_1 CB@13_mAd415_2 CB@13_mAd416_1 CB@13_mAd416_2 CB@13_mAd417_1 
+CB@13_mAd417_2 CB@13_mAd420_1 CB@13_mAd420_2 CB@13_mAd421_1 CB@13_mAd421_2 CB@13_mAd422_1 CB@13_mAd422_2 CB@13_mAd423_1 CB@13_mAd423_2 CB@13_mAd424_1 CB@13_mAd424_2 CB@13_mAd425_1 CB@13_mAd425_2 CB@13_mAd426_1 CB@13_mAd426_2 CB@13_mAd427_1 CB@13_mAd427_2 CB@13_mAd430_1 CB@13_mAd430_2 CB@13_mAd431_1 CB@13_mAd431_2 CB@13_mAd432_1 CB@13_mAd432_2 CB@13_mAd433_1 CB@13_mAd433_2 CB@13_mAd434_1 CB@13_mAd434_2 CB@13_mAd435_1 CB@13_mAd435_2 CB@13_mAd436_1 CB@13_mAd436_2 CB@13_mAd437_1 CB@13_mAd437_2 CB@13_mAd440_1 
+CB@13_mAd440_2 CB@13_mAd441_1 CB@13_mAd441_2 CB@13_mAd442_1 CB@13_mAd442_2 CB@13_mAd443_1 CB@13_mAd443_2 CB@13_mAd444_1 CB@13_mAd444_2 CB@13_mAd445_1 CB@13_mAd445_2 CB@13_mAd446_1 CB@13_mAd446_2 CB@13_mAd447_1 CB@13_mAd447_2 CB@13_mAd450_1 CB@13_mAd450_2 CB@13_mAd451_1 CB@13_mAd451_2 CB@13_mAd452_1 CB@13_mAd452_2 CB@13_mAd453_1 CB@13_mAd453_2 CB@13_mAd454_1 CB@13_mAd454_2 CB@13_mAd455_1 CB@13_mAd455_2 CB@13_mAd456_1 CB@13_mAd456_2 CB@13_mAd457_1 CB@13_mAd457_2 CB@13_mAd460_1 CB@13_mAd460_2 CB@13_mAd466_1 
+CB@13_mAd466_2 CB@13_mAd467_1 CB@13_mAd467_2 CB@13_mAd500_1 CB@13_mAd500_2 CB@13_mAd501_1 CB@13_mAd501_2 CB@13_mAd502_1 CB@13_mAd502_2 CB@13_mAd508_1 CB@13_mAd508_2 CB@13_mAd509_1 CB@13_mAd509_2 CB@13_mAd512_1 CB@13_mAd512_2 CB@13_mAd513_1 CB@13_mAd513_2 CB@13_mAd514_1 CB@13_mAd514_2 CB@13_mAd515_1 CB@13_mAd515_2 CB@13_mAd516_1 CB@13_mAd516_2 CB@13_mAd517_1 CB@13_mAd517_2 CB@13_mAd520_1 CB@13_mAd520_2 CB@13_mAd521_1 CB@13_mAd521_2 CB@13_mAd522_1 CB@13_mAd522_2 CB@13_mAd523_1 CB@13_mAd523_2 CB@13_mAd524_1 
+CB@13_mAd524_2 CB@13_mAd525_1 CB@13_mAd525_2 CB@13_mAd526_1 CB@13_mAd526_2 CB@13_mAd527_1 CB@13_mAd527_2 CB@13_mAd530_1 CB@13_mAd530_2 CB@13_mAd531_1 CB@13_mAd531_2 CB@13_mAd532_1 CB@13_mAd532_2 CB@13_mAd533_1 CB@13_mAd533_2 CB@13_mAd534_1 CB@13_mAd534_2 CB@13_mAd535_1 CB@13_mAd535_2 CB@13_mAd536_1 CB@13_mAd536_2 CB@13_mAd537_1 CB@13_mAd537_2 CB@13_mAd540_1 CB@13_mAd540_2 CB@13_mAd541_1 CB@13_mAd541_2 CB@13_mAd542_1 CB@13_mAd542_2 CB@13_mAd543_1 CB@13_mAd543_2 CB@13_mAd544_1 CB@13_mAd544_2 CB@13_mAd545_1 
+CB@13_mAd545_2 CB@13_mAd546_1 CB@13_mAd546_2 CB@13_mAd547_1 CB@13_mAd547_2 CB@13_mAd550_1 CB@13_mAd550_2 CB@13_mAd551_1 CB@13_mAd551_2 CB@13_mAd552_1 CB@13_mAd552_2 CB@13_mAd553_1 CB@13_mAd553_2 CB@13_mAd554_1 CB@13_mAd554_2 CB@13_mAd555_1 CB@13_mAd555_2 CB@13_mAd556_1 CB@13_mAd556_2 CB@13_mAd557_1 CB@13_mAd557_2 CB@13_mAd560_1 CB@13_mAd560_2 CB@13_mAd561_1 CB@13_mAd561_2 CB@13_mAd562_1 CB@13_mAd562_2 CB@13_mAd563_1 CB@13_mAd563_2 CB@13_mAd564_1 CB@13_mAd564_2 CB@13_mAd565_1 CB@13_mAd565_2 CB@13_mAd566_1 
+CB@13_mAd566_2 CB@13_mAd567_1 CB@13_mAd567_2 CB@13_mAd570_1 CB@13_mAd570_2 CB@13_mAd571_1 CB@13_mAd571_2 CB@13_mAd572_1 CB@13_mAd572_2 CB@13_mAd573_1 CB@13_mAd573_2 CB@13_mAd575_1 CB@13_mAd575_2 CB@13_mAd576_1 CB@13_mAd576_2 CB@13_mAd577_1 CB@13_mAd577_2 CB@13_mAd600_1 CB@13_mAd600_2 CB@13_mAd601_1 CB@13_mAd601_2 CB@13_mAd602_1 CB@13_mAd602_2 CB@13_mAd604_1 CB@13_mAd604_2 CB@13_mAd605_1 CB@13_mAd605_2 CB@13_mAd606_1 CB@13_mAd606_2 CB@13_mAd607_1 CB@13_mAd607_2 CB@13_mAd610_1 CB@13_mAd610_2 CB@13_mAd611_1 
+CB@13_mAd611_2 CB@13_mAd612_1 CB@13_mAd612_2 CB@13_mAd613_1 CB@13_mAd613_2 CB@13_mAd614_1 CB@13_mAd614_2 CB@13_mAd615_1 CB@13_mAd615_2 CB@13_mAd616_1 CB@13_mAd616_2 CB@13_mAd617_1 CB@13_mAd617_2 CB@13_mAd620_1 CB@13_mAd620_2 CB@13_mAd621_1 CB@13_mAd621_2 CB@13_mAd622_1 CB@13_mAd622_2 CB@13_mAd623_1 CB@13_mAd623_2 CB@13_mAd624_1 CB@13_mAd624_2 CB@13_mAd625_1 CB@13_mAd625_2 CB@13_mAd626_1 CB@13_mAd626_2 CB@13_mAd627_1 CB@13_mAd627_2 CB@13_mAd630_1 CB@13_mAd630_2 CB@13_mAd631_1 CB@13_mAd631_2 CB@13_mAd632_1 
+CB@13_mAd632_2 CB@13_mAd633_1 CB@13_mAd633_2 CB@13_mAd634_1 CB@13_mAd634_2 CB@13_mAd635_1 CB@13_mAd635_2 CB@13_mAd636_1 CB@13_mAd636_2 CB@13_mAd637_1 CB@13_mAd637_2 CB@13_mAd640_1 CB@13_mAd640_2 CB@13_mAd641_1 CB@13_mAd641_2 CB@13_mAd642_1 CB@13_mAd642_2 CB@13_mAd643_1 CB@13_mAd643_2 CB@13_mAd644_1 CB@13_mAd644_2 CB@13_mAd645_1 CB@13_mAd645_2 CB@13_mAd646_1 CB@13_mAd646_2 CB@13_mAd647_1 CB@13_mAd647_2 CB@13_mAd650_1 CB@13_mAd650_2 CB@13_mAd651_1 CB@13_mAd651_2 CB@13_mAd652_1 CB@13_mAd652_2 CB@13_mAd653_1 
+CB@13_mAd653_2 CB@13_mAd654_1 CB@13_mAd654_2 CB@13_mAd655_1 CB@13_mAd655_2 CB@13_mAd656_1 CB@13_mAd656_2 CB@13_mAd657_1 CB@13_mAd657_2 CB@13_mAd660_1 CB@13_mAd660_2 CB@13_mAd661_1 CB@13_mAd661_2 CB@13_mAd662_1 CB@13_mAd662_2 CB@13_mAd663_1 CB@13_mAd663_2 CB@13_mAd664_1 CB@13_mAd664_2 CB@13_mAd665_1 CB@13_mAd665_2 CB@13_mAd666_1 CB@13_mAd666_2 CB@13_mAd667_1 CB@13_mAd667_2 CB@13_mAd675_1 CB@13_mAd675_2 CB@13_mAd676_1 CB@13_mAd676_2 CB@13_mAd677_1 CB@13_mAd677_2 CB@13_mAd700_1 CB@13_mAd700_2 CB@13_mAd710_1 
+CB@13_mAd710_2 CB@13_mAd711_1 CB@13_mAd711_2 CB@13_mAd717_1 CB@13_mAd717_2 CB@13_mAd720_1 CB@13_mAd720_2 CB@13_mAd721_1 CB@13_mAd721_2 CB@13_mAd722_1 CB@13_mAd722_2 CB@13_mAd723_1 CB@13_mAd723_2 CB@13_mAd724_1 CB@13_mAd724_2 CB@13_mAd725_1 CB@13_mAd725_2 CB@13_mAd726_1 CB@13_mAd726_2 CB@13_mAd727_1 CB@13_mAd727_2 CB@13_mAd730_1 CB@13_mAd730_2 CB@13_mAd731_1 CB@13_mAd731_2 CB@13_mAd732_1 CB@13_mAd732_2 CB@13_mAd733_1 CB@13_mAd733_2 CB@13_mAd734_1 CB@13_mAd734_2 CB@13_mAd735_1 CB@13_mAd735_2 CB@13_mAd736_1 
+CB@13_mAd736_2 CB@13_mAd737_1 CB@13_mAd737_2 CB@13_mAd740_1 CB@13_mAd740_2 CB@13_mAd741_1 CB@13_mAd741_2 CB@13_mAd742_1 CB@13_mAd742_2 CB@13_mAd743_1 CB@13_mAd743_2 CB@13_mAd744_1 CB@13_mAd744_2 CB@13_mAd745_1 CB@13_mAd745_2 CB@13_mAd746_1 CB@13_mAd746_2 CB@13_mAd747_1 CB@13_mAd747_2 CB@13_mAd750_1 CB@13_mAd750_2 CB@13_mAd751_1 CB@13_mAd751_2 CB@13_mAd752_1 CB@13_mAd752_2 CB@13_mAd753_1 CB@13_mAd753_2 CB@13_mAd754_1 CB@13_mAd754_2 CB@13_mAd755_1 CB@13_mAd755_2 CB@13_mAd756_1 CB@13_mAd756_2 CB@13_mAd757_1 
+CB@13_mAd757_2 CB@13_mAd760_1 CB@13_mAd760_2 CB@13_mAd761_1 CB@13_mAd761_2 CB@13_mAd762_1 CB@13_mAd762_2 CB@13_mAd763_1 CB@13_mAd763_2 CB@13_mAd764_1 CB@13_mAd764_2 CB@13_mAd765_1 CB@13_mAd765_2 CB@13_mAd766_1 CB@13_mAd766_2 CB@13_mAd767_1 CB@13_mAd767_2 CB@13_mAd771_1 CB@13_mAd771_2 CB@13_mAd772_1 CB@13_mAd772_2 CB@13_mAd773_1 CB@13_mAd773_2 CB@13_mAd774_1 CB@13_mAd774_2 CB@13_mAd775_1 CB@13_mAd775_2 CB@13_mAd776_1 CB@13_mAd776_2 CB@13_mAd777_1 CB@13_mAd777_2 CB@13_X0 CB@13_X1 CB@13_X10 CB@13_X11 
+CB@13_X12 CB@13_X13 CB@13_X2 CB@13_X3 CB@13_X4 CB@13_X5 CB@13_X6 CB@13_X7 CB@13_X8 CB@13_X9 CB@13_Y1 CB@13_Y10 CB@13_Y11 CB@13_Y12 CB@13_Y2 CB@13_Y3 CB@13_Y4 CB@13_Y5 CB@13_Y6 CB@13_Y7 CB@13_Y8 CB@13_Y9 CB@13_Z1 CB@13_Z10 CB@13_Z11 CB@13_Z12 CB@13_Z2 CB@13_Z3 CB@13_Z4 CB@13_Z5 CB@13_Z6 CB@13_Z7 CB@13_Z8 CB@13_Z9 _5400TP094__CB
XCB@14 CB@14_K0 CB@14_K1 CB@14_K10 CB@14_K11 CB@14_K12 CB@14_K13 CB@14_K2 CB@14_K3 CB@14_K4 CB@14_K5 CB@14_K6 CB@14_K7 CB@14_K8 CB@14_K9 CB@14_mAd000_1 CB@14_mAd000_2 CB@14_mAd001_1 CB@14_mAd001_2 CB@14_mAd002_1 CB@14_mAd002_2 CB@14_mAd003_1 CB@14_mAd003_2 CB@14_mAd004_1 CB@14_mAd004_2 CB@14_mAd005_1 CB@14_mAd005_2 CB@14_mAd006_1 CB@14_mAd006_2 CB@14_mAd007_1 CB@14_mAd007_2 CB@14_mAd010_1 CB@14_mAd010_2 CB@14_mAd011_1 CB@14_mAd011_2 CB@14_mAd012_1 CB@14_mAd012_2 CB@14_mAd013_1 CB@14_mAd013_2 CB@14_mAd014_1 
+CB@14_mAd014_2 CB@14_mAd015_1 CB@14_mAd015_2 CB@14_mAd016_1 CB@14_mAd016_2 CB@14_mAd017_1 CB@14_mAd017_2 CB@14_mAd020_1 CB@14_mAd020_2 CB@14_mAd021_1 CB@14_mAd021_2 CB@14_mAd022_1 CB@14_mAd022_2 CB@14_mAd023_1 CB@14_mAd023_2 CB@14_mAd024_1 CB@14_mAd024_2 CB@14_mAd025_1 CB@14_mAd025_2 CB@14_mAd026_1 CB@14_mAd026_2 CB@14_mAd027_1 CB@14_mAd027_2 CB@14_mAd030_1 CB@14_mAd030_2 CB@14_mAd031_1 CB@14_mAd031_2 CB@14_mAd032_1 CB@14_mAd032_2 CB@14_mAd033_1 CB@14_mAd033_2 CB@14_mAd034_1 CB@14_mAd034_2 CB@14_mAd035_1 
+CB@14_mAd035_2 CB@14_mAd036_1 CB@14_mAd036_2 CB@14_mAd037_1 CB@14_mAd037_2 CB@14_mAd040_1 CB@14_mAd040_2 CB@14_mAd041_1 CB@14_mAd041_2 CB@14_mAd042_1 CB@14_mAd042_2 CB@14_mAd043_1 CB@14_mAd043_2 CB@14_mAd044_1 CB@14_mAd044_2 CB@14_mAd045_1 CB@14_mAd045_2 CB@14_mAd046_1 CB@14_mAd046_2 CB@14_mAd047_1 CB@14_mAd047_2 CB@14_mAd050_1 CB@14_mAd050_2 CB@14_mAd051_1 CB@14_mAd051_2 CB@14_mAd052_1 CB@14_mAd052_2 CB@14_mAd053_1 CB@14_mAd053_2 CB@14_mAd054_1 CB@14_mAd054_2 CB@14_mAd055_1 CB@14_mAd055_2 CB@14_mAd056_1 
+CB@14_mAd056_2 CB@14_mAd057_1 CB@14_mAd057_2 CB@14_mAd060_1 CB@14_mAd060_2 CB@14_mAd066_1 CB@14_mAd066_2 CB@14_mAd067_1 CB@14_mAd067_2 CB@14_mAd100_1 CB@14_mAd100_2 CB@14_mAd101_1 CB@14_mAd101_2 CB@14_mAd102_1 CB@14_mAd102_2 CB@14_mAd110_1 CB@14_mAd110_2 CB@14_mAd111_1 CB@14_mAd111_2 CB@14_mAd112_1 CB@14_mAd112_2 CB@14_mAd113_1 CB@14_mAd113_2 CB@14_mAd114_1 CB@14_mAd114_2 CB@14_mAd115_1 CB@14_mAd115_2 CB@14_mAd116_1 CB@14_mAd116_2 CB@14_mAd117_1 CB@14_mAd117_2 CB@14_mAd120_1 CB@14_mAd120_2 CB@14_mAd121_1 
+CB@14_mAd121_2 CB@14_mAd122_1 CB@14_mAd122_2 CB@14_mAd123_1 CB@14_mAd123_2 CB@14_mAd124_1 CB@14_mAd124_2 CB@14_mAd125_1 CB@14_mAd125_2 CB@14_mAd126_1 CB@14_mAd126_2 CB@14_mAd127_1 CB@14_mAd127_2 CB@14_mAd130_1 CB@14_mAd130_2 CB@14_mAd131_1 CB@14_mAd131_2 CB@14_mAd132_1 CB@14_mAd132_2 CB@14_mAd133_1 CB@14_mAd133_2 CB@14_mAd134_1 CB@14_mAd134_2 CB@14_mAd135_1 CB@14_mAd135_2 CB@14_mAd136_1 CB@14_mAd136_2 CB@14_mAd137_1 CB@14_mAd137_2 CB@14_mAd140_1 CB@14_mAd140_2 CB@14_mAd141_1 CB@14_mAd141_2 CB@14_mAd142_1 
+CB@14_mAd142_2 CB@14_mAd143_1 CB@14_mAd143_2 CB@14_mAd144_1 CB@14_mAd144_2 CB@14_mAd145_1 CB@14_mAd145_2 CB@14_mAd146_1 CB@14_mAd146_2 CB@14_mAd147_1 CB@14_mAd147_2 CB@14_mAd150_1 CB@14_mAd150_2 CB@14_mAd151_1 CB@14_mAd151_2 CB@14_mAd152_1 CB@14_mAd152_2 CB@14_mAd153_1 CB@14_mAd153_2 CB@14_mAd154_1 CB@14_mAd154_2 CB@14_mAd155_1 CB@14_mAd155_2 CB@14_mAd156_1 CB@14_mAd156_2 CB@14_mAd157_1 CB@14_mAd157_2 CB@14_mAd160_1 CB@14_mAd160_2 CB@14_mAd161_1 CB@14_mAd161_2 CB@14_mAd162_1 CB@14_mAd162_2 CB@14_mAd163_1 
+CB@14_mAd163_2 CB@14_mAd164_1 CB@14_mAd164_2 CB@14_mAd165_1 CB@14_mAd165_2 CB@14_mAd166_1 CB@14_mAd166_2 CB@14_mAd167_1 CB@14_mAd167_2 CB@14_mAd170_1 CB@14_mAd170_2 CB@14_mAd171_1 CB@14_mAd171_2 CB@14_mAd172_1 CB@14_mAd172_2 CB@14_mAd173_1 CB@14_mAd173_2 CB@14_mAd175_1 CB@14_mAd175_2 CB@14_mAd176_1 CB@14_mAd176_2 CB@14_mAd177_1 CB@14_mAd177_2 CB@14_mAd200_1 CB@14_mAd200_2 CB@14_mAd201_1 CB@14_mAd201_2 CB@14_mAd202_1 CB@14_mAd202_2 CB@14_mAd204_1 CB@14_mAd204_2 CB@14_mAd205_1 CB@14_mAd205_2 CB@14_mAd206_1 
+CB@14_mAd206_2 CB@14_mAd207_1 CB@14_mAd207_2 CB@14_mAd210_1 CB@14_mAd210_2 CB@14_mAd211_1 CB@14_mAd211_2 CB@14_mAd212_1 CB@14_mAd212_2 CB@14_mAd213_1 CB@14_mAd213_2 CB@14_mAd214_1 CB@14_mAd214_2 CB@14_mAd215_1 CB@14_mAd215_2 CB@14_mAd216_1 CB@14_mAd216_2 CB@14_mAd217_1 CB@14_mAd217_2 CB@14_mAd220_1 CB@14_mAd220_2 CB@14_mAd221_1 CB@14_mAd221_2 CB@14_mAd222_1 CB@14_mAd222_2 CB@14_mAd223_1 CB@14_mAd223_2 CB@14_mAd224_1 CB@14_mAd224_2 CB@14_mAd225_1 CB@14_mAd225_2 CB@14_mAd226_1 CB@14_mAd226_2 CB@14_mAd227_1 
+CB@14_mAd227_2 CB@14_mAd230_1 CB@14_mAd230_2 CB@14_mAd231_1 CB@14_mAd231_2 CB@14_mAd232_1 CB@14_mAd232_2 CB@14_mAd233_1 CB@14_mAd233_2 CB@14_mAd234_1 CB@14_mAd234_2 CB@14_mAd235_1 CB@14_mAd235_2 CB@14_mAd236_1 CB@14_mAd236_2 CB@14_mAd237_1 CB@14_mAd237_2 CB@14_mAd240_1 CB@14_mAd240_2 CB@14_mAd241_1 CB@14_mAd241_2 CB@14_mAd242_1 CB@14_mAd242_2 CB@14_mAd243_1 CB@14_mAd243_2 CB@14_mAd244_1 CB@14_mAd244_2 CB@14_mAd245_1 CB@14_mAd245_2 CB@14_mAd246_1 CB@14_mAd246_2 CB@14_mAd247_1 CB@14_mAd247_2 CB@14_mAd250_1 
+CB@14_mAd250_2 CB@14_mAd251_1 CB@14_mAd251_2 CB@14_mAd252_1 CB@14_mAd252_2 CB@14_mAd253_1 CB@14_mAd253_2 CB@14_mAd254_1 CB@14_mAd254_2 CB@14_mAd255_1 CB@14_mAd255_2 CB@14_mAd256_1 CB@14_mAd256_2 CB@14_mAd257_1 CB@14_mAd257_2 CB@14_mAd260_1 CB@14_mAd260_2 CB@14_mAd261_1 CB@14_mAd261_2 CB@14_mAd262_1 CB@14_mAd262_2 CB@14_mAd263_1 CB@14_mAd263_2 CB@14_mAd264_1 CB@14_mAd264_2 CB@14_mAd265_1 CB@14_mAd265_2 CB@14_mAd266_1 CB@14_mAd266_2 CB@14_mAd267_1 CB@14_mAd267_2 CB@14_mAd275_1 CB@14_mAd275_2 CB@14_mAd276_1 
+CB@14_mAd276_2 CB@14_mAd277_1 CB@14_mAd277_2 CB@14_mAd300_1 CB@14_mAd300_2 CB@14_mAd310_1 CB@14_mAd310_2 CB@14_mAd311_1 CB@14_mAd311_2 CB@14_mAd317_1 CB@14_mAd317_2 CB@14_mAd320_1 CB@14_mAd320_2 CB@14_mAd321_1 CB@14_mAd321_2 CB@14_mAd322_1 CB@14_mAd322_2 CB@14_mAd323_1 CB@14_mAd323_2 CB@14_mAd324_1 CB@14_mAd324_2 CB@14_mAd325_1 CB@14_mAd325_2 CB@14_mAd326_1 CB@14_mAd326_2 CB@14_mAd327_1 CB@14_mAd327_2 CB@14_mAd330_1 CB@14_mAd330_2 CB@14_mAd331_1 CB@14_mAd331_2 CB@14_mAd332_1 CB@14_mAd332_2 CB@14_mAd333_1 
+CB@14_mAd333_2 CB@14_mAd334_1 CB@14_mAd334_2 CB@14_mAd335_1 CB@14_mAd335_2 CB@14_mAd336_1 CB@14_mAd336_2 CB@14_mAd337_1 CB@14_mAd337_2 CB@14_mAd340_1 CB@14_mAd340_2 CB@14_mAd341_1 CB@14_mAd341_2 CB@14_mAd342_1 CB@14_mAd342_2 CB@14_mAd343_1 CB@14_mAd343_2 CB@14_mAd344_1 CB@14_mAd344_2 CB@14_mAd345_1 CB@14_mAd345_2 CB@14_mAd346_1 CB@14_mAd346_2 CB@14_mAd347_1 CB@14_mAd347_2 CB@14_mAd350_1 CB@14_mAd350_2 CB@14_mAd351_1 CB@14_mAd351_2 CB@14_mAd352_1 CB@14_mAd352_2 CB@14_mAd353_1 CB@14_mAd353_2 CB@14_mAd354_1 
+CB@14_mAd354_2 CB@14_mAd355_1 CB@14_mAd355_2 CB@14_mAd356_1 CB@14_mAd356_2 CB@14_mAd357_1 CB@14_mAd357_2 CB@14_mAd360_1 CB@14_mAd360_2 CB@14_mAd361_1 CB@14_mAd361_2 CB@14_mAd362_1 CB@14_mAd362_2 CB@14_mAd363_1 CB@14_mAd363_2 CB@14_mAd364_1 CB@14_mAd364_2 CB@14_mAd365_1 CB@14_mAd365_2 CB@14_mAd366_1 CB@14_mAd366_2 CB@14_mAd367_1 CB@14_mAd367_2 CB@14_mAd371_1 CB@14_mAd371_2 CB@14_mAd372_1 CB@14_mAd372_2 CB@14_mAd373_1 CB@14_mAd373_2 CB@14_mAd374_1 CB@14_mAd374_2 CB@14_mAd375_1 CB@14_mAd375_2 CB@14_mAd376_1 
+CB@14_mAd376_2 CB@14_mAd377_1 CB@14_mAd377_2 CB@14_mAd400_1 CB@14_mAd400_2 CB@14_mAd401_1 CB@14_mAd401_2 CB@14_mAd402_1 CB@14_mAd402_2 CB@14_mAd403_1 CB@14_mAd403_2 CB@14_mAd404_1 CB@14_mAd404_2 CB@14_mAd405_1 CB@14_mAd405_2 CB@14_mAd406_1 CB@14_mAd406_2 CB@14_mAd407_1 CB@14_mAd407_2 CB@14_mAd410_1 CB@14_mAd410_2 CB@14_mAd411_1 CB@14_mAd411_2 CB@14_mAd412_1 CB@14_mAd412_2 CB@14_mAd413_1 CB@14_mAd413_2 CB@14_mAd414_1 CB@14_mAd414_2 CB@14_mAd415_1 CB@14_mAd415_2 CB@14_mAd416_1 CB@14_mAd416_2 CB@14_mAd417_1 
+CB@14_mAd417_2 CB@14_mAd420_1 CB@14_mAd420_2 CB@14_mAd421_1 CB@14_mAd421_2 CB@14_mAd422_1 CB@14_mAd422_2 CB@14_mAd423_1 CB@14_mAd423_2 CB@14_mAd424_1 CB@14_mAd424_2 CB@14_mAd425_1 CB@14_mAd425_2 CB@14_mAd426_1 CB@14_mAd426_2 CB@14_mAd427_1 CB@14_mAd427_2 CB@14_mAd430_1 CB@14_mAd430_2 CB@14_mAd431_1 CB@14_mAd431_2 CB@14_mAd432_1 CB@14_mAd432_2 CB@14_mAd433_1 CB@14_mAd433_2 CB@14_mAd434_1 CB@14_mAd434_2 CB@14_mAd435_1 CB@14_mAd435_2 CB@14_mAd436_1 CB@14_mAd436_2 CB@14_mAd437_1 CB@14_mAd437_2 CB@14_mAd440_1 
+CB@14_mAd440_2 CB@14_mAd441_1 CB@14_mAd441_2 CB@14_mAd442_1 CB@14_mAd442_2 CB@14_mAd443_1 CB@14_mAd443_2 CB@14_mAd444_1 CB@14_mAd444_2 CB@14_mAd445_1 CB@14_mAd445_2 CB@14_mAd446_1 CB@14_mAd446_2 CB@14_mAd447_1 CB@14_mAd447_2 CB@14_mAd450_1 CB@14_mAd450_2 CB@14_mAd451_1 CB@14_mAd451_2 CB@14_mAd452_1 CB@14_mAd452_2 CB@14_mAd453_1 CB@14_mAd453_2 CB@14_mAd454_1 CB@14_mAd454_2 CB@14_mAd455_1 CB@14_mAd455_2 CB@14_mAd456_1 CB@14_mAd456_2 CB@14_mAd457_1 CB@14_mAd457_2 CB@14_mAd460_1 CB@14_mAd460_2 CB@14_mAd466_1 
+CB@14_mAd466_2 CB@14_mAd467_1 CB@14_mAd467_2 CB@14_mAd500_1 CB@14_mAd500_2 CB@14_mAd501_1 CB@14_mAd501_2 CB@14_mAd502_1 CB@14_mAd502_2 CB@14_mAd508_1 CB@14_mAd508_2 CB@14_mAd509_1 CB@14_mAd509_2 CB@14_mAd512_1 CB@14_mAd512_2 CB@14_mAd513_1 CB@14_mAd513_2 CB@14_mAd514_1 CB@14_mAd514_2 CB@14_mAd515_1 CB@14_mAd515_2 CB@14_mAd516_1 CB@14_mAd516_2 CB@14_mAd517_1 CB@14_mAd517_2 CB@14_mAd520_1 CB@14_mAd520_2 CB@14_mAd521_1 CB@14_mAd521_2 CB@14_mAd522_1 CB@14_mAd522_2 CB@14_mAd523_1 CB@14_mAd523_2 CB@14_mAd524_1 
+CB@14_mAd524_2 CB@14_mAd525_1 CB@14_mAd525_2 CB@14_mAd526_1 CB@14_mAd526_2 CB@14_mAd527_1 CB@14_mAd527_2 CB@14_mAd530_1 CB@14_mAd530_2 CB@14_mAd531_1 CB@14_mAd531_2 CB@14_mAd532_1 CB@14_mAd532_2 CB@14_mAd533_1 CB@14_mAd533_2 CB@14_mAd534_1 CB@14_mAd534_2 CB@14_mAd535_1 CB@14_mAd535_2 CB@14_mAd536_1 CB@14_mAd536_2 CB@14_mAd537_1 CB@14_mAd537_2 CB@14_mAd540_1 CB@14_mAd540_2 CB@14_mAd541_1 CB@14_mAd541_2 CB@14_mAd542_1 CB@14_mAd542_2 CB@14_mAd543_1 CB@14_mAd543_2 CB@14_mAd544_1 CB@14_mAd544_2 CB@14_mAd545_1 
+CB@14_mAd545_2 CB@14_mAd546_1 CB@14_mAd546_2 CB@14_mAd547_1 CB@14_mAd547_2 CB@14_mAd550_1 CB@14_mAd550_2 CB@14_mAd551_1 CB@14_mAd551_2 CB@14_mAd552_1 CB@14_mAd552_2 CB@14_mAd553_1 CB@14_mAd553_2 CB@14_mAd554_1 CB@14_mAd554_2 CB@14_mAd555_1 CB@14_mAd555_2 CB@14_mAd556_1 CB@14_mAd556_2 CB@14_mAd557_1 CB@14_mAd557_2 CB@14_mAd560_1 CB@14_mAd560_2 CB@14_mAd561_1 CB@14_mAd561_2 CB@14_mAd562_1 CB@14_mAd562_2 CB@14_mAd563_1 CB@14_mAd563_2 CB@14_mAd564_1 CB@14_mAd564_2 CB@14_mAd565_1 CB@14_mAd565_2 CB@14_mAd566_1 
+CB@14_mAd566_2 CB@14_mAd567_1 CB@14_mAd567_2 CB@14_mAd570_1 CB@14_mAd570_2 CB@14_mAd571_1 CB@14_mAd571_2 CB@14_mAd572_1 CB@14_mAd572_2 CB@14_mAd573_1 CB@14_mAd573_2 CB@14_mAd575_1 CB@14_mAd575_2 CB@14_mAd576_1 CB@14_mAd576_2 CB@14_mAd577_1 CB@14_mAd577_2 CB@14_mAd600_1 CB@14_mAd600_2 CB@14_mAd601_1 CB@14_mAd601_2 CB@14_mAd602_1 CB@14_mAd602_2 CB@14_mAd604_1 CB@14_mAd604_2 CB@14_mAd605_1 CB@14_mAd605_2 CB@14_mAd606_1 CB@14_mAd606_2 CB@14_mAd607_1 CB@14_mAd607_2 CB@14_mAd610_1 CB@14_mAd610_2 CB@14_mAd611_1 
+CB@14_mAd611_2 CB@14_mAd612_1 CB@14_mAd612_2 CB@14_mAd613_1 CB@14_mAd613_2 CB@14_mAd614_1 CB@14_mAd614_2 CB@14_mAd615_1 CB@14_mAd615_2 CB@14_mAd616_1 CB@14_mAd616_2 CB@14_mAd617_1 CB@14_mAd617_2 CB@14_mAd620_1 CB@14_mAd620_2 CB@14_mAd621_1 CB@14_mAd621_2 CB@14_mAd622_1 CB@14_mAd622_2 CB@14_mAd623_1 CB@14_mAd623_2 CB@14_mAd624_1 CB@14_mAd624_2 CB@14_mAd625_1 CB@14_mAd625_2 CB@14_mAd626_1 CB@14_mAd626_2 CB@14_mAd627_1 CB@14_mAd627_2 CB@14_mAd630_1 CB@14_mAd630_2 CB@14_mAd631_1 CB@14_mAd631_2 CB@14_mAd632_1 
+CB@14_mAd632_2 CB@14_mAd633_1 CB@14_mAd633_2 CB@14_mAd634_1 CB@14_mAd634_2 CB@14_mAd635_1 CB@14_mAd635_2 CB@14_mAd636_1 CB@14_mAd636_2 CB@14_mAd637_1 CB@14_mAd637_2 CB@14_mAd640_1 CB@14_mAd640_2 CB@14_mAd641_1 CB@14_mAd641_2 CB@14_mAd642_1 CB@14_mAd642_2 CB@14_mAd643_1 CB@14_mAd643_2 CB@14_mAd644_1 CB@14_mAd644_2 CB@14_mAd645_1 CB@14_mAd645_2 CB@14_mAd646_1 CB@14_mAd646_2 CB@14_mAd647_1 CB@14_mAd647_2 CB@14_mAd650_1 CB@14_mAd650_2 CB@14_mAd651_1 CB@14_mAd651_2 CB@14_mAd652_1 CB@14_mAd652_2 CB@14_mAd653_1 
+CB@14_mAd653_2 CB@14_mAd654_1 CB@14_mAd654_2 CB@14_mAd655_1 CB@14_mAd655_2 CB@14_mAd656_1 CB@14_mAd656_2 CB@14_mAd657_1 CB@14_mAd657_2 CB@14_mAd660_1 CB@14_mAd660_2 CB@14_mAd661_1 CB@14_mAd661_2 CB@14_mAd662_1 CB@14_mAd662_2 CB@14_mAd663_1 CB@14_mAd663_2 CB@14_mAd664_1 CB@14_mAd664_2 CB@14_mAd665_1 CB@14_mAd665_2 CB@14_mAd666_1 CB@14_mAd666_2 CB@14_mAd667_1 CB@14_mAd667_2 CB@14_mAd675_1 CB@14_mAd675_2 CB@14_mAd676_1 CB@14_mAd676_2 CB@14_mAd677_1 CB@14_mAd677_2 CB@14_mAd700_1 CB@14_mAd700_2 CB@14_mAd710_1 
+CB@14_mAd710_2 CB@14_mAd711_1 CB@14_mAd711_2 CB@14_mAd717_1 CB@14_mAd717_2 CB@14_mAd720_1 CB@14_mAd720_2 CB@14_mAd721_1 CB@14_mAd721_2 CB@14_mAd722_1 CB@14_mAd722_2 CB@14_mAd723_1 CB@14_mAd723_2 CB@14_mAd724_1 CB@14_mAd724_2 CB@14_mAd725_1 CB@14_mAd725_2 CB@14_mAd726_1 CB@14_mAd726_2 CB@14_mAd727_1 CB@14_mAd727_2 CB@14_mAd730_1 CB@14_mAd730_2 CB@14_mAd731_1 CB@14_mAd731_2 CB@14_mAd732_1 CB@14_mAd732_2 CB@14_mAd733_1 CB@14_mAd733_2 CB@14_mAd734_1 CB@14_mAd734_2 CB@14_mAd735_1 CB@14_mAd735_2 CB@14_mAd736_1 
+CB@14_mAd736_2 CB@14_mAd737_1 CB@14_mAd737_2 CB@14_mAd740_1 CB@14_mAd740_2 CB@14_mAd741_1 CB@14_mAd741_2 CB@14_mAd742_1 CB@14_mAd742_2 CB@14_mAd743_1 CB@14_mAd743_2 CB@14_mAd744_1 CB@14_mAd744_2 CB@14_mAd745_1 CB@14_mAd745_2 CB@14_mAd746_1 CB@14_mAd746_2 CB@14_mAd747_1 CB@14_mAd747_2 CB@14_mAd750_1 CB@14_mAd750_2 CB@14_mAd751_1 CB@14_mAd751_2 CB@14_mAd752_1 CB@14_mAd752_2 CB@14_mAd753_1 CB@14_mAd753_2 CB@14_mAd754_1 CB@14_mAd754_2 CB@14_mAd755_1 CB@14_mAd755_2 CB@14_mAd756_1 CB@14_mAd756_2 CB@14_mAd757_1 
+CB@14_mAd757_2 CB@14_mAd760_1 CB@14_mAd760_2 CB@14_mAd761_1 CB@14_mAd761_2 CB@14_mAd762_1 CB@14_mAd762_2 CB@14_mAd763_1 CB@14_mAd763_2 CB@14_mAd764_1 CB@14_mAd764_2 CB@14_mAd765_1 CB@14_mAd765_2 CB@14_mAd766_1 CB@14_mAd766_2 CB@14_mAd767_1 CB@14_mAd767_2 CB@14_mAd771_1 CB@14_mAd771_2 CB@14_mAd772_1 CB@14_mAd772_2 CB@14_mAd773_1 CB@14_mAd773_2 CB@14_mAd774_1 CB@14_mAd774_2 CB@14_mAd775_1 CB@14_mAd775_2 CB@14_mAd776_1 CB@14_mAd776_2 CB@14_mAd777_1 CB@14_mAd777_2 CB@14_X0 CB@14_X1 CB@14_X10 CB@14_X11 
+CB@14_X12 CB@14_X13 CB@14_X2 CB@14_X3 CB@14_X4 CB@14_X5 CB@14_X6 CB@14_X7 CB@14_X8 CB@14_X9 CB@14_Y1 CB@14_Y10 CB@14_Y11 CB@14_Y12 CB@14_Y2 CB@14_Y3 CB@14_Y4 CB@14_Y5 CB@14_Y6 CB@14_Y7 CB@14_Y8 CB@14_Y9 CB@14_Z1 CB@14_Z10 CB@14_Z11 CB@14_Z12 CB@14_Z2 CB@14_Z3 CB@14_Z4 CB@14_Z5 CB@14_Z6 CB@14_Z7 CB@14_Z8 CB@14_Z9 _5400TP094__CB
XCB@15 CB@15_K0 CB@15_K1 CB@15_K10 CB@15_K11 CB@15_K12 CB@15_K13 CB@15_K2 CB@15_K3 CB@15_K4 CB@15_K5 CB@15_K6 CB@15_K7 CB@15_K8 CB@15_K9 CB@15_mAd000_1 CB@15_mAd000_2 CB@15_mAd001_1 CB@15_mAd001_2 CB@15_mAd002_1 CB@15_mAd002_2 CB@15_mAd003_1 CB@15_mAd003_2 CB@15_mAd004_1 CB@15_mAd004_2 CB@15_mAd005_1 CB@15_mAd005_2 CB@15_mAd006_1 CB@15_mAd006_2 CB@15_mAd007_1 CB@15_mAd007_2 CB@15_mAd010_1 CB@15_mAd010_2 CB@15_mAd011_1 CB@15_mAd011_2 CB@15_mAd012_1 CB@15_mAd012_2 CB@15_mAd013_1 CB@15_mAd013_2 CB@15_mAd014_1 
+CB@15_mAd014_2 CB@15_mAd015_1 CB@15_mAd015_2 CB@15_mAd016_1 CB@15_mAd016_2 CB@15_mAd017_1 CB@15_mAd017_2 CB@15_mAd020_1 CB@15_mAd020_2 CB@15_mAd021_1 CB@15_mAd021_2 CB@15_mAd022_1 CB@15_mAd022_2 CB@15_mAd023_1 CB@15_mAd023_2 CB@15_mAd024_1 CB@15_mAd024_2 CB@15_mAd025_1 CB@15_mAd025_2 CB@15_mAd026_1 CB@15_mAd026_2 CB@15_mAd027_1 CB@15_mAd027_2 CB@15_mAd030_1 CB@15_mAd030_2 CB@15_mAd031_1 CB@15_mAd031_2 CB@15_mAd032_1 CB@15_mAd032_2 CB@15_mAd033_1 CB@15_mAd033_2 CB@15_mAd034_1 CB@15_mAd034_2 CB@15_mAd035_1 
+CB@15_mAd035_2 CB@15_mAd036_1 CB@15_mAd036_2 CB@15_mAd037_1 CB@15_mAd037_2 CB@15_mAd040_1 CB@15_mAd040_2 CB@15_mAd041_1 CB@15_mAd041_2 CB@15_mAd042_1 CB@15_mAd042_2 CB@15_mAd043_1 CB@15_mAd043_2 CB@15_mAd044_1 CB@15_mAd044_2 CB@15_mAd045_1 CB@15_mAd045_2 CB@15_mAd046_1 CB@15_mAd046_2 CB@15_mAd047_1 CB@15_mAd047_2 CB@15_mAd050_1 CB@15_mAd050_2 CB@15_mAd051_1 CB@15_mAd051_2 CB@15_mAd052_1 CB@15_mAd052_2 CB@15_mAd053_1 CB@15_mAd053_2 CB@15_mAd054_1 CB@15_mAd054_2 CB@15_mAd055_1 CB@15_mAd055_2 CB@15_mAd056_1 
+CB@15_mAd056_2 CB@15_mAd057_1 CB@15_mAd057_2 CB@15_mAd060_1 CB@15_mAd060_2 CB@15_mAd066_1 CB@15_mAd066_2 CB@15_mAd067_1 CB@15_mAd067_2 CB@15_mAd100_1 CB@15_mAd100_2 CB@15_mAd101_1 CB@15_mAd101_2 CB@15_mAd102_1 CB@15_mAd102_2 CB@15_mAd110_1 CB@15_mAd110_2 CB@15_mAd111_1 CB@15_mAd111_2 CB@15_mAd112_1 CB@15_mAd112_2 CB@15_mAd113_1 CB@15_mAd113_2 CB@15_mAd114_1 CB@15_mAd114_2 CB@15_mAd115_1 CB@15_mAd115_2 CB@15_mAd116_1 CB@15_mAd116_2 CB@15_mAd117_1 CB@15_mAd117_2 CB@15_mAd120_1 CB@15_mAd120_2 CB@15_mAd121_1 
+CB@15_mAd121_2 CB@15_mAd122_1 CB@15_mAd122_2 CB@15_mAd123_1 CB@15_mAd123_2 CB@15_mAd124_1 CB@15_mAd124_2 CB@15_mAd125_1 CB@15_mAd125_2 CB@15_mAd126_1 CB@15_mAd126_2 CB@15_mAd127_1 CB@15_mAd127_2 CB@15_mAd130_1 CB@15_mAd130_2 CB@15_mAd131_1 CB@15_mAd131_2 CB@15_mAd132_1 CB@15_mAd132_2 CB@15_mAd133_1 CB@15_mAd133_2 CB@15_mAd134_1 CB@15_mAd134_2 CB@15_mAd135_1 CB@15_mAd135_2 CB@15_mAd136_1 CB@15_mAd136_2 CB@15_mAd137_1 CB@15_mAd137_2 CB@15_mAd140_1 CB@15_mAd140_2 CB@15_mAd141_1 CB@15_mAd141_2 CB@15_mAd142_1 
+CB@15_mAd142_2 CB@15_mAd143_1 CB@15_mAd143_2 CB@15_mAd144_1 CB@15_mAd144_2 CB@15_mAd145_1 CB@15_mAd145_2 CB@15_mAd146_1 CB@15_mAd146_2 CB@15_mAd147_1 CB@15_mAd147_2 CB@15_mAd150_1 CB@15_mAd150_2 CB@15_mAd151_1 CB@15_mAd151_2 CB@15_mAd152_1 CB@15_mAd152_2 CB@15_mAd153_1 CB@15_mAd153_2 CB@15_mAd154_1 CB@15_mAd154_2 CB@15_mAd155_1 CB@15_mAd155_2 CB@15_mAd156_1 CB@15_mAd156_2 CB@15_mAd157_1 CB@15_mAd157_2 CB@15_mAd160_1 CB@15_mAd160_2 CB@15_mAd161_1 CB@15_mAd161_2 CB@15_mAd162_1 CB@15_mAd162_2 CB@15_mAd163_1 
+CB@15_mAd163_2 CB@15_mAd164_1 CB@15_mAd164_2 CB@15_mAd165_1 CB@15_mAd165_2 CB@15_mAd166_1 CB@15_mAd166_2 CB@15_mAd167_1 CB@15_mAd167_2 CB@15_mAd170_1 CB@15_mAd170_2 CB@15_mAd171_1 CB@15_mAd171_2 CB@15_mAd172_1 CB@15_mAd172_2 CB@15_mAd173_1 CB@15_mAd173_2 CB@15_mAd175_1 CB@15_mAd175_2 CB@15_mAd176_1 CB@15_mAd176_2 CB@15_mAd177_1 CB@15_mAd177_2 CB@15_mAd200_1 CB@15_mAd200_2 CB@15_mAd201_1 CB@15_mAd201_2 CB@15_mAd202_1 CB@15_mAd202_2 CB@15_mAd204_1 CB@15_mAd204_2 CB@15_mAd205_1 CB@15_mAd205_2 CB@15_mAd206_1 
+CB@15_mAd206_2 CB@15_mAd207_1 CB@15_mAd207_2 CB@15_mAd210_1 CB@15_mAd210_2 CB@15_mAd211_1 CB@15_mAd211_2 CB@15_mAd212_1 CB@15_mAd212_2 CB@15_mAd213_1 CB@15_mAd213_2 CB@15_mAd214_1 CB@15_mAd214_2 CB@15_mAd215_1 CB@15_mAd215_2 CB@15_mAd216_1 CB@15_mAd216_2 CB@15_mAd217_1 CB@15_mAd217_2 CB@15_mAd220_1 CB@15_mAd220_2 CB@15_mAd221_1 CB@15_mAd221_2 CB@15_mAd222_1 CB@15_mAd222_2 CB@15_mAd223_1 CB@15_mAd223_2 CB@15_mAd224_1 CB@15_mAd224_2 CB@15_mAd225_1 CB@15_mAd225_2 CB@15_mAd226_1 CB@15_mAd226_2 CB@15_mAd227_1 
+CB@15_mAd227_2 CB@15_mAd230_1 CB@15_mAd230_2 CB@15_mAd231_1 CB@15_mAd231_2 CB@15_mAd232_1 CB@15_mAd232_2 CB@15_mAd233_1 CB@15_mAd233_2 CB@15_mAd234_1 CB@15_mAd234_2 CB@15_mAd235_1 CB@15_mAd235_2 CB@15_mAd236_1 CB@15_mAd236_2 CB@15_mAd237_1 CB@15_mAd237_2 CB@15_mAd240_1 CB@15_mAd240_2 CB@15_mAd241_1 CB@15_mAd241_2 CB@15_mAd242_1 CB@15_mAd242_2 CB@15_mAd243_1 CB@15_mAd243_2 CB@15_mAd244_1 CB@15_mAd244_2 CB@15_mAd245_1 CB@15_mAd245_2 CB@15_mAd246_1 CB@15_mAd246_2 CB@15_mAd247_1 CB@15_mAd247_2 CB@15_mAd250_1 
+CB@15_mAd250_2 CB@15_mAd251_1 CB@15_mAd251_2 CB@15_mAd252_1 CB@15_mAd252_2 CB@15_mAd253_1 CB@15_mAd253_2 CB@15_mAd254_1 CB@15_mAd254_2 CB@15_mAd255_1 CB@15_mAd255_2 CB@15_mAd256_1 CB@15_mAd256_2 CB@15_mAd257_1 CB@15_mAd257_2 CB@15_mAd260_1 CB@15_mAd260_2 CB@15_mAd261_1 CB@15_mAd261_2 CB@15_mAd262_1 CB@15_mAd262_2 CB@15_mAd263_1 CB@15_mAd263_2 CB@15_mAd264_1 CB@15_mAd264_2 CB@15_mAd265_1 CB@15_mAd265_2 CB@15_mAd266_1 CB@15_mAd266_2 CB@15_mAd267_1 CB@15_mAd267_2 CB@15_mAd275_1 CB@15_mAd275_2 CB@15_mAd276_1 
+CB@15_mAd276_2 CB@15_mAd277_1 CB@15_mAd277_2 CB@15_mAd300_1 CB@15_mAd300_2 CB@15_mAd310_1 CB@15_mAd310_2 CB@15_mAd311_1 CB@15_mAd311_2 CB@15_mAd317_1 CB@15_mAd317_2 CB@15_mAd320_1 CB@15_mAd320_2 CB@15_mAd321_1 CB@15_mAd321_2 CB@15_mAd322_1 CB@15_mAd322_2 CB@15_mAd323_1 CB@15_mAd323_2 CB@15_mAd324_1 CB@15_mAd324_2 CB@15_mAd325_1 CB@15_mAd325_2 CB@15_mAd326_1 CB@15_mAd326_2 CB@15_mAd327_1 CB@15_mAd327_2 CB@15_mAd330_1 CB@15_mAd330_2 CB@15_mAd331_1 CB@15_mAd331_2 CB@15_mAd332_1 CB@15_mAd332_2 CB@15_mAd333_1 
+CB@15_mAd333_2 CB@15_mAd334_1 CB@15_mAd334_2 CB@15_mAd335_1 CB@15_mAd335_2 CB@15_mAd336_1 CB@15_mAd336_2 CB@15_mAd337_1 CB@15_mAd337_2 CB@15_mAd340_1 CB@15_mAd340_2 CB@15_mAd341_1 CB@15_mAd341_2 CB@15_mAd342_1 CB@15_mAd342_2 CB@15_mAd343_1 CB@15_mAd343_2 CB@15_mAd344_1 CB@15_mAd344_2 CB@15_mAd345_1 CB@15_mAd345_2 CB@15_mAd346_1 CB@15_mAd346_2 CB@15_mAd347_1 CB@15_mAd347_2 CB@15_mAd350_1 CB@15_mAd350_2 CB@15_mAd351_1 CB@15_mAd351_2 CB@15_mAd352_1 CB@15_mAd352_2 CB@15_mAd353_1 CB@15_mAd353_2 CB@15_mAd354_1 
+CB@15_mAd354_2 CB@15_mAd355_1 CB@15_mAd355_2 CB@15_mAd356_1 CB@15_mAd356_2 CB@15_mAd357_1 CB@15_mAd357_2 CB@15_mAd360_1 CB@15_mAd360_2 CB@15_mAd361_1 CB@15_mAd361_2 CB@15_mAd362_1 CB@15_mAd362_2 CB@15_mAd363_1 CB@15_mAd363_2 CB@15_mAd364_1 CB@15_mAd364_2 CB@15_mAd365_1 CB@15_mAd365_2 CB@15_mAd366_1 CB@15_mAd366_2 CB@15_mAd367_1 CB@15_mAd367_2 CB@15_mAd371_1 CB@15_mAd371_2 CB@15_mAd372_1 CB@15_mAd372_2 CB@15_mAd373_1 CB@15_mAd373_2 CB@15_mAd374_1 CB@15_mAd374_2 CB@15_mAd375_1 CB@15_mAd375_2 CB@15_mAd376_1 
+CB@15_mAd376_2 CB@15_mAd377_1 CB@15_mAd377_2 CB@15_mAd400_1 CB@15_mAd400_2 CB@15_mAd401_1 CB@15_mAd401_2 CB@15_mAd402_1 CB@15_mAd402_2 CB@15_mAd403_1 CB@15_mAd403_2 CB@15_mAd404_1 CB@15_mAd404_2 CB@15_mAd405_1 CB@15_mAd405_2 CB@15_mAd406_1 CB@15_mAd406_2 CB@15_mAd407_1 CB@15_mAd407_2 CB@15_mAd410_1 CB@15_mAd410_2 CB@15_mAd411_1 CB@15_mAd411_2 CB@15_mAd412_1 CB@15_mAd412_2 CB@15_mAd413_1 CB@15_mAd413_2 CB@15_mAd414_1 CB@15_mAd414_2 CB@15_mAd415_1 CB@15_mAd415_2 CB@15_mAd416_1 CB@15_mAd416_2 CB@15_mAd417_1 
+CB@15_mAd417_2 CB@15_mAd420_1 CB@15_mAd420_2 CB@15_mAd421_1 CB@15_mAd421_2 CB@15_mAd422_1 CB@15_mAd422_2 CB@15_mAd423_1 CB@15_mAd423_2 CB@15_mAd424_1 CB@15_mAd424_2 CB@15_mAd425_1 CB@15_mAd425_2 CB@15_mAd426_1 CB@15_mAd426_2 CB@15_mAd427_1 CB@15_mAd427_2 CB@15_mAd430_1 CB@15_mAd430_2 CB@15_mAd431_1 CB@15_mAd431_2 CB@15_mAd432_1 CB@15_mAd432_2 CB@15_mAd433_1 CB@15_mAd433_2 CB@15_mAd434_1 CB@15_mAd434_2 CB@15_mAd435_1 CB@15_mAd435_2 CB@15_mAd436_1 CB@15_mAd436_2 CB@15_mAd437_1 CB@15_mAd437_2 CB@15_mAd440_1 
+CB@15_mAd440_2 CB@15_mAd441_1 CB@15_mAd441_2 CB@15_mAd442_1 CB@15_mAd442_2 CB@15_mAd443_1 CB@15_mAd443_2 CB@15_mAd444_1 CB@15_mAd444_2 CB@15_mAd445_1 CB@15_mAd445_2 CB@15_mAd446_1 CB@15_mAd446_2 CB@15_mAd447_1 CB@15_mAd447_2 CB@15_mAd450_1 CB@15_mAd450_2 CB@15_mAd451_1 CB@15_mAd451_2 CB@15_mAd452_1 CB@15_mAd452_2 CB@15_mAd453_1 CB@15_mAd453_2 CB@15_mAd454_1 CB@15_mAd454_2 CB@15_mAd455_1 CB@15_mAd455_2 CB@15_mAd456_1 CB@15_mAd456_2 CB@15_mAd457_1 CB@15_mAd457_2 CB@15_mAd460_1 CB@15_mAd460_2 CB@15_mAd466_1 
+CB@15_mAd466_2 CB@15_mAd467_1 CB@15_mAd467_2 CB@15_mAd500_1 CB@15_mAd500_2 CB@15_mAd501_1 CB@15_mAd501_2 CB@15_mAd502_1 CB@15_mAd502_2 CB@15_mAd508_1 CB@15_mAd508_2 CB@15_mAd509_1 CB@15_mAd509_2 CB@15_mAd512_1 CB@15_mAd512_2 CB@15_mAd513_1 CB@15_mAd513_2 CB@15_mAd514_1 CB@15_mAd514_2 CB@15_mAd515_1 CB@15_mAd515_2 CB@15_mAd516_1 CB@15_mAd516_2 CB@15_mAd517_1 CB@15_mAd517_2 CB@15_mAd520_1 CB@15_mAd520_2 CB@15_mAd521_1 CB@15_mAd521_2 CB@15_mAd522_1 CB@15_mAd522_2 CB@15_mAd523_1 CB@15_mAd523_2 CB@15_mAd524_1 
+CB@15_mAd524_2 CB@15_mAd525_1 CB@15_mAd525_2 CB@15_mAd526_1 CB@15_mAd526_2 CB@15_mAd527_1 CB@15_mAd527_2 CB@15_mAd530_1 CB@15_mAd530_2 CB@15_mAd531_1 CB@15_mAd531_2 CB@15_mAd532_1 CB@15_mAd532_2 CB@15_mAd533_1 CB@15_mAd533_2 CB@15_mAd534_1 CB@15_mAd534_2 CB@15_mAd535_1 CB@15_mAd535_2 CB@15_mAd536_1 CB@15_mAd536_2 CB@15_mAd537_1 CB@15_mAd537_2 CB@15_mAd540_1 CB@15_mAd540_2 CB@15_mAd541_1 CB@15_mAd541_2 CB@15_mAd542_1 CB@15_mAd542_2 CB@15_mAd543_1 CB@15_mAd543_2 CB@15_mAd544_1 CB@15_mAd544_2 CB@15_mAd545_1 
+CB@15_mAd545_2 CB@15_mAd546_1 CB@15_mAd546_2 CB@15_mAd547_1 CB@15_mAd547_2 CB@15_mAd550_1 CB@15_mAd550_2 CB@15_mAd551_1 CB@15_mAd551_2 CB@15_mAd552_1 CB@15_mAd552_2 CB@15_mAd553_1 CB@15_mAd553_2 CB@15_mAd554_1 CB@15_mAd554_2 CB@15_mAd555_1 CB@15_mAd555_2 CB@15_mAd556_1 CB@15_mAd556_2 CB@15_mAd557_1 CB@15_mAd557_2 CB@15_mAd560_1 CB@15_mAd560_2 CB@15_mAd561_1 CB@15_mAd561_2 CB@15_mAd562_1 CB@15_mAd562_2 CB@15_mAd563_1 CB@15_mAd563_2 CB@15_mAd564_1 CB@15_mAd564_2 CB@15_mAd565_1 CB@15_mAd565_2 CB@15_mAd566_1 
+CB@15_mAd566_2 CB@15_mAd567_1 CB@15_mAd567_2 CB@15_mAd570_1 CB@15_mAd570_2 CB@15_mAd571_1 CB@15_mAd571_2 CB@15_mAd572_1 CB@15_mAd572_2 CB@15_mAd573_1 CB@15_mAd573_2 CB@15_mAd575_1 CB@15_mAd575_2 CB@15_mAd576_1 CB@15_mAd576_2 CB@15_mAd577_1 CB@15_mAd577_2 CB@15_mAd600_1 CB@15_mAd600_2 CB@15_mAd601_1 CB@15_mAd601_2 CB@15_mAd602_1 CB@15_mAd602_2 CB@15_mAd604_1 CB@15_mAd604_2 CB@15_mAd605_1 CB@15_mAd605_2 CB@15_mAd606_1 CB@15_mAd606_2 CB@15_mAd607_1 CB@15_mAd607_2 CB@15_mAd610_1 CB@15_mAd610_2 CB@15_mAd611_1 
+CB@15_mAd611_2 CB@15_mAd612_1 CB@15_mAd612_2 CB@15_mAd613_1 CB@15_mAd613_2 CB@15_mAd614_1 CB@15_mAd614_2 CB@15_mAd615_1 CB@15_mAd615_2 CB@15_mAd616_1 CB@15_mAd616_2 CB@15_mAd617_1 CB@15_mAd617_2 CB@15_mAd620_1 CB@15_mAd620_2 CB@15_mAd621_1 CB@15_mAd621_2 CB@15_mAd622_1 CB@15_mAd622_2 CB@15_mAd623_1 CB@15_mAd623_2 CB@15_mAd624_1 CB@15_mAd624_2 CB@15_mAd625_1 CB@15_mAd625_2 CB@15_mAd626_1 CB@15_mAd626_2 CB@15_mAd627_1 CB@15_mAd627_2 CB@15_mAd630_1 CB@15_mAd630_2 CB@15_mAd631_1 CB@15_mAd631_2 CB@15_mAd632_1 
+CB@15_mAd632_2 CB@15_mAd633_1 CB@15_mAd633_2 CB@15_mAd634_1 CB@15_mAd634_2 CB@15_mAd635_1 CB@15_mAd635_2 CB@15_mAd636_1 CB@15_mAd636_2 CB@15_mAd637_1 CB@15_mAd637_2 CB@15_mAd640_1 CB@15_mAd640_2 CB@15_mAd641_1 CB@15_mAd641_2 CB@15_mAd642_1 CB@15_mAd642_2 CB@15_mAd643_1 CB@15_mAd643_2 CB@15_mAd644_1 CB@15_mAd644_2 CB@15_mAd645_1 CB@15_mAd645_2 CB@15_mAd646_1 CB@15_mAd646_2 CB@15_mAd647_1 CB@15_mAd647_2 CB@15_mAd650_1 CB@15_mAd650_2 CB@15_mAd651_1 CB@15_mAd651_2 CB@15_mAd652_1 CB@15_mAd652_2 CB@15_mAd653_1 
+CB@15_mAd653_2 CB@15_mAd654_1 CB@15_mAd654_2 CB@15_mAd655_1 CB@15_mAd655_2 CB@15_mAd656_1 CB@15_mAd656_2 CB@15_mAd657_1 CB@15_mAd657_2 CB@15_mAd660_1 CB@15_mAd660_2 CB@15_mAd661_1 CB@15_mAd661_2 CB@15_mAd662_1 CB@15_mAd662_2 CB@15_mAd663_1 CB@15_mAd663_2 CB@15_mAd664_1 CB@15_mAd664_2 CB@15_mAd665_1 CB@15_mAd665_2 CB@15_mAd666_1 CB@15_mAd666_2 CB@15_mAd667_1 CB@15_mAd667_2 CB@15_mAd675_1 CB@15_mAd675_2 CB@15_mAd676_1 CB@15_mAd676_2 CB@15_mAd677_1 CB@15_mAd677_2 CB@15_mAd700_1 CB@15_mAd700_2 CB@15_mAd710_1 
+CB@15_mAd710_2 CB@15_mAd711_1 CB@15_mAd711_2 CB@15_mAd717_1 CB@15_mAd717_2 CB@15_mAd720_1 CB@15_mAd720_2 CB@15_mAd721_1 CB@15_mAd721_2 CB@15_mAd722_1 CB@15_mAd722_2 CB@15_mAd723_1 CB@15_mAd723_2 CB@15_mAd724_1 CB@15_mAd724_2 CB@15_mAd725_1 CB@15_mAd725_2 CB@15_mAd726_1 CB@15_mAd726_2 CB@15_mAd727_1 CB@15_mAd727_2 CB@15_mAd730_1 CB@15_mAd730_2 CB@15_mAd731_1 CB@15_mAd731_2 CB@15_mAd732_1 CB@15_mAd732_2 CB@15_mAd733_1 CB@15_mAd733_2 CB@15_mAd734_1 CB@15_mAd734_2 CB@15_mAd735_1 CB@15_mAd735_2 CB@15_mAd736_1 
+CB@15_mAd736_2 CB@15_mAd737_1 CB@15_mAd737_2 CB@15_mAd740_1 CB@15_mAd740_2 CB@15_mAd741_1 CB@15_mAd741_2 CB@15_mAd742_1 CB@15_mAd742_2 CB@15_mAd743_1 CB@15_mAd743_2 CB@15_mAd744_1 CB@15_mAd744_2 CB@15_mAd745_1 CB@15_mAd745_2 CB@15_mAd746_1 CB@15_mAd746_2 CB@15_mAd747_1 CB@15_mAd747_2 CB@15_mAd750_1 CB@15_mAd750_2 CB@15_mAd751_1 CB@15_mAd751_2 CB@15_mAd752_1 CB@15_mAd752_2 CB@15_mAd753_1 CB@15_mAd753_2 CB@15_mAd754_1 CB@15_mAd754_2 CB@15_mAd755_1 CB@15_mAd755_2 CB@15_mAd756_1 CB@15_mAd756_2 CB@15_mAd757_1 
+CB@15_mAd757_2 CB@15_mAd760_1 CB@15_mAd760_2 CB@15_mAd761_1 CB@15_mAd761_2 CB@15_mAd762_1 CB@15_mAd762_2 CB@15_mAd763_1 CB@15_mAd763_2 CB@15_mAd764_1 CB@15_mAd764_2 CB@15_mAd765_1 CB@15_mAd765_2 CB@15_mAd766_1 CB@15_mAd766_2 CB@15_mAd767_1 CB@15_mAd767_2 CB@15_mAd771_1 CB@15_mAd771_2 CB@15_mAd772_1 CB@15_mAd772_2 CB@15_mAd773_1 CB@15_mAd773_2 CB@15_mAd774_1 CB@15_mAd774_2 CB@15_mAd775_1 CB@15_mAd775_2 CB@15_mAd776_1 CB@15_mAd776_2 CB@15_mAd777_1 CB@15_mAd777_2 CB@15_X0 CB@15_X1 CB@15_X10 CB@15_X11 
+CB@15_X12 CB@15_X13 CB@15_X2 CB@15_X3 CB@15_X4 CB@15_X5 CB@15_X6 CB@15_X7 CB@15_X8 CB@15_X9 CB@15_Y1 CB@15_Y10 CB@15_Y11 CB@15_Y12 CB@15_Y2 CB@15_Y3 CB@15_Y4 CB@15_Y5 CB@15_Y6 CB@15_Y7 CB@15_Y8 CB@15_Y9 CB@15_Z1 CB@15_Z10 CB@15_Z11 CB@15_Z12 CB@15_Z2 CB@15_Z3 CB@15_Z4 CB@15_Z5 CB@15_Z6 CB@15_Z7 CB@15_Z8 CB@15_Z9 _5400TP094__CB
XCB@16 CB@16_K0 CB@16_K1 CB@16_K10 CB@16_K11 CB@16_K12 CB@16_K13 CB@16_K2 CB@16_K3 CB@16_K4 CB@16_K5 CB@16_K6 CB@16_K7 CB@16_K8 CB@16_K9 CB@16_mAd000_1 CB@16_mAd000_2 CB@16_mAd001_1 CB@16_mAd001_2 CB@16_mAd002_1 CB@16_mAd002_2 CB@16_mAd003_1 CB@16_mAd003_2 CB@16_mAd004_1 CB@16_mAd004_2 CB@16_mAd005_1 CB@16_mAd005_2 CB@16_mAd006_1 CB@16_mAd006_2 CB@16_mAd007_1 CB@16_mAd007_2 CB@16_mAd010_1 CB@16_mAd010_2 CB@16_mAd011_1 CB@16_mAd011_2 CB@16_mAd012_1 CB@16_mAd012_2 CB@16_mAd013_1 CB@16_mAd013_2 CB@16_mAd014_1 
+CB@16_mAd014_2 CB@16_mAd015_1 CB@16_mAd015_2 CB@16_mAd016_1 CB@16_mAd016_2 CB@16_mAd017_1 CB@16_mAd017_2 CB@16_mAd020_1 CB@16_mAd020_2 CB@16_mAd021_1 CB@16_mAd021_2 CB@16_mAd022_1 CB@16_mAd022_2 CB@16_mAd023_1 CB@16_mAd023_2 CB@16_mAd024_1 CB@16_mAd024_2 CB@16_mAd025_1 CB@16_mAd025_2 CB@16_mAd026_1 CB@16_mAd026_2 CB@16_mAd027_1 CB@16_mAd027_2 CB@16_mAd030_1 CB@16_mAd030_2 CB@16_mAd031_1 CB@16_mAd031_2 CB@16_mAd032_1 CB@16_mAd032_2 CB@16_mAd033_1 CB@16_mAd033_2 CB@16_mAd034_1 CB@16_mAd034_2 CB@16_mAd035_1 
+CB@16_mAd035_2 CB@16_mAd036_1 CB@16_mAd036_2 CB@16_mAd037_1 CB@16_mAd037_2 CB@16_mAd040_1 CB@16_mAd040_2 CB@16_mAd041_1 CB@16_mAd041_2 CB@16_mAd042_1 CB@16_mAd042_2 CB@16_mAd043_1 CB@16_mAd043_2 CB@16_mAd044_1 CB@16_mAd044_2 CB@16_mAd045_1 CB@16_mAd045_2 CB@16_mAd046_1 CB@16_mAd046_2 CB@16_mAd047_1 CB@16_mAd047_2 CB@16_mAd050_1 CB@16_mAd050_2 CB@16_mAd051_1 CB@16_mAd051_2 CB@16_mAd052_1 CB@16_mAd052_2 CB@16_mAd053_1 CB@16_mAd053_2 CB@16_mAd054_1 CB@16_mAd054_2 CB@16_mAd055_1 CB@16_mAd055_2 CB@16_mAd056_1 
+CB@16_mAd056_2 CB@16_mAd057_1 CB@16_mAd057_2 CB@16_mAd060_1 CB@16_mAd060_2 CB@16_mAd066_1 CB@16_mAd066_2 CB@16_mAd067_1 CB@16_mAd067_2 CB@16_mAd100_1 CB@16_mAd100_2 CB@16_mAd101_1 CB@16_mAd101_2 CB@16_mAd102_1 CB@16_mAd102_2 CB@16_mAd110_1 CB@16_mAd110_2 CB@16_mAd111_1 CB@16_mAd111_2 CB@16_mAd112_1 CB@16_mAd112_2 CB@16_mAd113_1 CB@16_mAd113_2 CB@16_mAd114_1 CB@16_mAd114_2 CB@16_mAd115_1 CB@16_mAd115_2 CB@16_mAd116_1 CB@16_mAd116_2 CB@16_mAd117_1 CB@16_mAd117_2 CB@16_mAd120_1 CB@16_mAd120_2 CB@16_mAd121_1 
+CB@16_mAd121_2 CB@16_mAd122_1 CB@16_mAd122_2 CB@16_mAd123_1 CB@16_mAd123_2 CB@16_mAd124_1 CB@16_mAd124_2 CB@16_mAd125_1 CB@16_mAd125_2 CB@16_mAd126_1 CB@16_mAd126_2 CB@16_mAd127_1 CB@16_mAd127_2 CB@16_mAd130_1 CB@16_mAd130_2 CB@16_mAd131_1 CB@16_mAd131_2 CB@16_mAd132_1 CB@16_mAd132_2 CB@16_mAd133_1 CB@16_mAd133_2 CB@16_mAd134_1 CB@16_mAd134_2 CB@16_mAd135_1 CB@16_mAd135_2 CB@16_mAd136_1 CB@16_mAd136_2 CB@16_mAd137_1 CB@16_mAd137_2 CB@16_mAd140_1 CB@16_mAd140_2 CB@16_mAd141_1 CB@16_mAd141_2 CB@16_mAd142_1 
+CB@16_mAd142_2 CB@16_mAd143_1 CB@16_mAd143_2 CB@16_mAd144_1 CB@16_mAd144_2 CB@16_mAd145_1 CB@16_mAd145_2 CB@16_mAd146_1 CB@16_mAd146_2 CB@16_mAd147_1 CB@16_mAd147_2 CB@16_mAd150_1 CB@16_mAd150_2 CB@16_mAd151_1 CB@16_mAd151_2 CB@16_mAd152_1 CB@16_mAd152_2 CB@16_mAd153_1 CB@16_mAd153_2 CB@16_mAd154_1 CB@16_mAd154_2 CB@16_mAd155_1 CB@16_mAd155_2 CB@16_mAd156_1 CB@16_mAd156_2 CB@16_mAd157_1 CB@16_mAd157_2 CB@16_mAd160_1 CB@16_mAd160_2 CB@16_mAd161_1 CB@16_mAd161_2 CB@16_mAd162_1 CB@16_mAd162_2 CB@16_mAd163_1 
+CB@16_mAd163_2 CB@16_mAd164_1 CB@16_mAd164_2 CB@16_mAd165_1 CB@16_mAd165_2 CB@16_mAd166_1 CB@16_mAd166_2 CB@16_mAd167_1 CB@16_mAd167_2 CB@16_mAd170_1 CB@16_mAd170_2 CB@16_mAd171_1 CB@16_mAd171_2 CB@16_mAd172_1 CB@16_mAd172_2 CB@16_mAd173_1 CB@16_mAd173_2 CB@16_mAd175_1 CB@16_mAd175_2 CB@16_mAd176_1 CB@16_mAd176_2 CB@16_mAd177_1 CB@16_mAd177_2 CB@16_mAd200_1 CB@16_mAd200_2 CB@16_mAd201_1 CB@16_mAd201_2 CB@16_mAd202_1 CB@16_mAd202_2 CB@16_mAd204_1 CB@16_mAd204_2 CB@16_mAd205_1 CB@16_mAd205_2 CB@16_mAd206_1 
+CB@16_mAd206_2 CB@16_mAd207_1 CB@16_mAd207_2 CB@16_mAd210_1 CB@16_mAd210_2 CB@16_mAd211_1 CB@16_mAd211_2 CB@16_mAd212_1 CB@16_mAd212_2 CB@16_mAd213_1 CB@16_mAd213_2 CB@16_mAd214_1 CB@16_mAd214_2 CB@16_mAd215_1 CB@16_mAd215_2 CB@16_mAd216_1 CB@16_mAd216_2 CB@16_mAd217_1 CB@16_mAd217_2 CB@16_mAd220_1 CB@16_mAd220_2 CB@16_mAd221_1 CB@16_mAd221_2 CB@16_mAd222_1 CB@16_mAd222_2 CB@16_mAd223_1 CB@16_mAd223_2 CB@16_mAd224_1 CB@16_mAd224_2 CB@16_mAd225_1 CB@16_mAd225_2 CB@16_mAd226_1 CB@16_mAd226_2 CB@16_mAd227_1 
+CB@16_mAd227_2 CB@16_mAd230_1 CB@16_mAd230_2 CB@16_mAd231_1 CB@16_mAd231_2 CB@16_mAd232_1 CB@16_mAd232_2 CB@16_mAd233_1 CB@16_mAd233_2 CB@16_mAd234_1 CB@16_mAd234_2 CB@16_mAd235_1 CB@16_mAd235_2 CB@16_mAd236_1 CB@16_mAd236_2 CB@16_mAd237_1 CB@16_mAd237_2 CB@16_mAd240_1 CB@16_mAd240_2 CB@16_mAd241_1 CB@16_mAd241_2 CB@16_mAd242_1 CB@16_mAd242_2 CB@16_mAd243_1 CB@16_mAd243_2 CB@16_mAd244_1 CB@16_mAd244_2 CB@16_mAd245_1 CB@16_mAd245_2 CB@16_mAd246_1 CB@16_mAd246_2 CB@16_mAd247_1 CB@16_mAd247_2 CB@16_mAd250_1 
+CB@16_mAd250_2 CB@16_mAd251_1 CB@16_mAd251_2 CB@16_mAd252_1 CB@16_mAd252_2 CB@16_mAd253_1 CB@16_mAd253_2 CB@16_mAd254_1 CB@16_mAd254_2 CB@16_mAd255_1 CB@16_mAd255_2 CB@16_mAd256_1 CB@16_mAd256_2 CB@16_mAd257_1 CB@16_mAd257_2 CB@16_mAd260_1 CB@16_mAd260_2 CB@16_mAd261_1 CB@16_mAd261_2 CB@16_mAd262_1 CB@16_mAd262_2 CB@16_mAd263_1 CB@16_mAd263_2 CB@16_mAd264_1 CB@16_mAd264_2 CB@16_mAd265_1 CB@16_mAd265_2 CB@16_mAd266_1 CB@16_mAd266_2 CB@16_mAd267_1 CB@16_mAd267_2 CB@16_mAd275_1 CB@16_mAd275_2 CB@16_mAd276_1 
+CB@16_mAd276_2 CB@16_mAd277_1 CB@16_mAd277_2 CB@16_mAd300_1 CB@16_mAd300_2 CB@16_mAd310_1 CB@16_mAd310_2 CB@16_mAd311_1 CB@16_mAd311_2 CB@16_mAd317_1 CB@16_mAd317_2 CB@16_mAd320_1 CB@16_mAd320_2 CB@16_mAd321_1 CB@16_mAd321_2 CB@16_mAd322_1 CB@16_mAd322_2 CB@16_mAd323_1 CB@16_mAd323_2 CB@16_mAd324_1 CB@16_mAd324_2 CB@16_mAd325_1 CB@16_mAd325_2 CB@16_mAd326_1 CB@16_mAd326_2 CB@16_mAd327_1 CB@16_mAd327_2 CB@16_mAd330_1 CB@16_mAd330_2 CB@16_mAd331_1 CB@16_mAd331_2 CB@16_mAd332_1 CB@16_mAd332_2 CB@16_mAd333_1 
+CB@16_mAd333_2 CB@16_mAd334_1 CB@16_mAd334_2 CB@16_mAd335_1 CB@16_mAd335_2 CB@16_mAd336_1 CB@16_mAd336_2 CB@16_mAd337_1 CB@16_mAd337_2 CB@16_mAd340_1 CB@16_mAd340_2 CB@16_mAd341_1 CB@16_mAd341_2 CB@16_mAd342_1 CB@16_mAd342_2 CB@16_mAd343_1 CB@16_mAd343_2 CB@16_mAd344_1 CB@16_mAd344_2 CB@16_mAd345_1 CB@16_mAd345_2 CB@16_mAd346_1 CB@16_mAd346_2 CB@16_mAd347_1 CB@16_mAd347_2 CB@16_mAd350_1 CB@16_mAd350_2 CB@16_mAd351_1 CB@16_mAd351_2 CB@16_mAd352_1 CB@16_mAd352_2 CB@16_mAd353_1 CB@16_mAd353_2 CB@16_mAd354_1 
+CB@16_mAd354_2 CB@16_mAd355_1 CB@16_mAd355_2 CB@16_mAd356_1 CB@16_mAd356_2 CB@16_mAd357_1 CB@16_mAd357_2 CB@16_mAd360_1 CB@16_mAd360_2 CB@16_mAd361_1 CB@16_mAd361_2 CB@16_mAd362_1 CB@16_mAd362_2 CB@16_mAd363_1 CB@16_mAd363_2 CB@16_mAd364_1 CB@16_mAd364_2 CB@16_mAd365_1 CB@16_mAd365_2 CB@16_mAd366_1 CB@16_mAd366_2 CB@16_mAd367_1 CB@16_mAd367_2 CB@16_mAd371_1 CB@16_mAd371_2 CB@16_mAd372_1 CB@16_mAd372_2 CB@16_mAd373_1 CB@16_mAd373_2 CB@16_mAd374_1 CB@16_mAd374_2 CB@16_mAd375_1 CB@16_mAd375_2 CB@16_mAd376_1 
+CB@16_mAd376_2 CB@16_mAd377_1 CB@16_mAd377_2 CB@16_mAd400_1 CB@16_mAd400_2 CB@16_mAd401_1 CB@16_mAd401_2 CB@16_mAd402_1 CB@16_mAd402_2 CB@16_mAd403_1 CB@16_mAd403_2 CB@16_mAd404_1 CB@16_mAd404_2 CB@16_mAd405_1 CB@16_mAd405_2 CB@16_mAd406_1 CB@16_mAd406_2 CB@16_mAd407_1 CB@16_mAd407_2 CB@16_mAd410_1 CB@16_mAd410_2 CB@16_mAd411_1 CB@16_mAd411_2 CB@16_mAd412_1 CB@16_mAd412_2 CB@16_mAd413_1 CB@16_mAd413_2 CB@16_mAd414_1 CB@16_mAd414_2 CB@16_mAd415_1 CB@16_mAd415_2 CB@16_mAd416_1 CB@16_mAd416_2 CB@16_mAd417_1 
+CB@16_mAd417_2 CB@16_mAd420_1 CB@16_mAd420_2 CB@16_mAd421_1 CB@16_mAd421_2 CB@16_mAd422_1 CB@16_mAd422_2 CB@16_mAd423_1 CB@16_mAd423_2 CB@16_mAd424_1 CB@16_mAd424_2 CB@16_mAd425_1 CB@16_mAd425_2 CB@16_mAd426_1 CB@16_mAd426_2 CB@16_mAd427_1 CB@16_mAd427_2 CB@16_mAd430_1 CB@16_mAd430_2 CB@16_mAd431_1 CB@16_mAd431_2 CB@16_mAd432_1 CB@16_mAd432_2 CB@16_mAd433_1 CB@16_mAd433_2 CB@16_mAd434_1 CB@16_mAd434_2 CB@16_mAd435_1 CB@16_mAd435_2 CB@16_mAd436_1 CB@16_mAd436_2 CB@16_mAd437_1 CB@16_mAd437_2 CB@16_mAd440_1 
+CB@16_mAd440_2 CB@16_mAd441_1 CB@16_mAd441_2 CB@16_mAd442_1 CB@16_mAd442_2 CB@16_mAd443_1 CB@16_mAd443_2 CB@16_mAd444_1 CB@16_mAd444_2 CB@16_mAd445_1 CB@16_mAd445_2 CB@16_mAd446_1 CB@16_mAd446_2 CB@16_mAd447_1 CB@16_mAd447_2 CB@16_mAd450_1 CB@16_mAd450_2 CB@16_mAd451_1 CB@16_mAd451_2 CB@16_mAd452_1 CB@16_mAd452_2 CB@16_mAd453_1 CB@16_mAd453_2 CB@16_mAd454_1 CB@16_mAd454_2 CB@16_mAd455_1 CB@16_mAd455_2 CB@16_mAd456_1 CB@16_mAd456_2 CB@16_mAd457_1 CB@16_mAd457_2 CB@16_mAd460_1 CB@16_mAd460_2 CB@16_mAd466_1 
+CB@16_mAd466_2 CB@16_mAd467_1 CB@16_mAd467_2 CB@16_mAd500_1 CB@16_mAd500_2 CB@16_mAd501_1 CB@16_mAd501_2 CB@16_mAd502_1 CB@16_mAd502_2 CB@16_mAd508_1 CB@16_mAd508_2 CB@16_mAd509_1 CB@16_mAd509_2 CB@16_mAd512_1 CB@16_mAd512_2 CB@16_mAd513_1 CB@16_mAd513_2 CB@16_mAd514_1 CB@16_mAd514_2 CB@16_mAd515_1 CB@16_mAd515_2 CB@16_mAd516_1 CB@16_mAd516_2 CB@16_mAd517_1 CB@16_mAd517_2 CB@16_mAd520_1 CB@16_mAd520_2 CB@16_mAd521_1 CB@16_mAd521_2 CB@16_mAd522_1 CB@16_mAd522_2 CB@16_mAd523_1 CB@16_mAd523_2 CB@16_mAd524_1 
+CB@16_mAd524_2 CB@16_mAd525_1 CB@16_mAd525_2 CB@16_mAd526_1 CB@16_mAd526_2 CB@16_mAd527_1 CB@16_mAd527_2 CB@16_mAd530_1 CB@16_mAd530_2 CB@16_mAd531_1 CB@16_mAd531_2 CB@16_mAd532_1 CB@16_mAd532_2 CB@16_mAd533_1 CB@16_mAd533_2 CB@16_mAd534_1 CB@16_mAd534_2 CB@16_mAd535_1 CB@16_mAd535_2 CB@16_mAd536_1 CB@16_mAd536_2 CB@16_mAd537_1 CB@16_mAd537_2 CB@16_mAd540_1 CB@16_mAd540_2 CB@16_mAd541_1 CB@16_mAd541_2 CB@16_mAd542_1 CB@16_mAd542_2 CB@16_mAd543_1 CB@16_mAd543_2 CB@16_mAd544_1 CB@16_mAd544_2 CB@16_mAd545_1 
+CB@16_mAd545_2 CB@16_mAd546_1 CB@16_mAd546_2 CB@16_mAd547_1 CB@16_mAd547_2 CB@16_mAd550_1 CB@16_mAd550_2 CB@16_mAd551_1 CB@16_mAd551_2 CB@16_mAd552_1 CB@16_mAd552_2 CB@16_mAd553_1 CB@16_mAd553_2 CB@16_mAd554_1 CB@16_mAd554_2 CB@16_mAd555_1 CB@16_mAd555_2 CB@16_mAd556_1 CB@16_mAd556_2 CB@16_mAd557_1 CB@16_mAd557_2 CB@16_mAd560_1 CB@16_mAd560_2 CB@16_mAd561_1 CB@16_mAd561_2 CB@16_mAd562_1 CB@16_mAd562_2 CB@16_mAd563_1 CB@16_mAd563_2 CB@16_mAd564_1 CB@16_mAd564_2 CB@16_mAd565_1 CB@16_mAd565_2 CB@16_mAd566_1 
+CB@16_mAd566_2 CB@16_mAd567_1 CB@16_mAd567_2 CB@16_mAd570_1 CB@16_mAd570_2 CB@16_mAd571_1 CB@16_mAd571_2 CB@16_mAd572_1 CB@16_mAd572_2 CB@16_mAd573_1 CB@16_mAd573_2 CB@16_mAd575_1 CB@16_mAd575_2 CB@16_mAd576_1 CB@16_mAd576_2 CB@16_mAd577_1 CB@16_mAd577_2 CB@16_mAd600_1 CB@16_mAd600_2 CB@16_mAd601_1 CB@16_mAd601_2 CB@16_mAd602_1 CB@16_mAd602_2 CB@16_mAd604_1 CB@16_mAd604_2 CB@16_mAd605_1 CB@16_mAd605_2 CB@16_mAd606_1 CB@16_mAd606_2 CB@16_mAd607_1 CB@16_mAd607_2 CB@16_mAd610_1 CB@16_mAd610_2 CB@16_mAd611_1 
+CB@16_mAd611_2 CB@16_mAd612_1 CB@16_mAd612_2 CB@16_mAd613_1 CB@16_mAd613_2 CB@16_mAd614_1 CB@16_mAd614_2 CB@16_mAd615_1 CB@16_mAd615_2 CB@16_mAd616_1 CB@16_mAd616_2 CB@16_mAd617_1 CB@16_mAd617_2 CB@16_mAd620_1 CB@16_mAd620_2 CB@16_mAd621_1 CB@16_mAd621_2 CB@16_mAd622_1 CB@16_mAd622_2 CB@16_mAd623_1 CB@16_mAd623_2 CB@16_mAd624_1 CB@16_mAd624_2 CB@16_mAd625_1 CB@16_mAd625_2 CB@16_mAd626_1 CB@16_mAd626_2 CB@16_mAd627_1 CB@16_mAd627_2 CB@16_mAd630_1 CB@16_mAd630_2 CB@16_mAd631_1 CB@16_mAd631_2 CB@16_mAd632_1 
+CB@16_mAd632_2 CB@16_mAd633_1 CB@16_mAd633_2 CB@16_mAd634_1 CB@16_mAd634_2 CB@16_mAd635_1 CB@16_mAd635_2 CB@16_mAd636_1 CB@16_mAd636_2 CB@16_mAd637_1 CB@16_mAd637_2 CB@16_mAd640_1 CB@16_mAd640_2 CB@16_mAd641_1 CB@16_mAd641_2 CB@16_mAd642_1 CB@16_mAd642_2 CB@16_mAd643_1 CB@16_mAd643_2 CB@16_mAd644_1 CB@16_mAd644_2 CB@16_mAd645_1 CB@16_mAd645_2 CB@16_mAd646_1 CB@16_mAd646_2 CB@16_mAd647_1 CB@16_mAd647_2 CB@16_mAd650_1 CB@16_mAd650_2 CB@16_mAd651_1 CB@16_mAd651_2 CB@16_mAd652_1 CB@16_mAd652_2 CB@16_mAd653_1 
+CB@16_mAd653_2 CB@16_mAd654_1 CB@16_mAd654_2 CB@16_mAd655_1 CB@16_mAd655_2 CB@16_mAd656_1 CB@16_mAd656_2 CB@16_mAd657_1 CB@16_mAd657_2 CB@16_mAd660_1 CB@16_mAd660_2 CB@16_mAd661_1 CB@16_mAd661_2 CB@16_mAd662_1 CB@16_mAd662_2 CB@16_mAd663_1 CB@16_mAd663_2 CB@16_mAd664_1 CB@16_mAd664_2 CB@16_mAd665_1 CB@16_mAd665_2 CB@16_mAd666_1 CB@16_mAd666_2 CB@16_mAd667_1 CB@16_mAd667_2 CB@16_mAd675_1 CB@16_mAd675_2 CB@16_mAd676_1 CB@16_mAd676_2 CB@16_mAd677_1 CB@16_mAd677_2 CB@16_mAd700_1 CB@16_mAd700_2 CB@16_mAd710_1 
+CB@16_mAd710_2 CB@16_mAd711_1 CB@16_mAd711_2 CB@16_mAd717_1 CB@16_mAd717_2 CB@16_mAd720_1 CB@16_mAd720_2 CB@16_mAd721_1 CB@16_mAd721_2 CB@16_mAd722_1 CB@16_mAd722_2 CB@16_mAd723_1 CB@16_mAd723_2 CB@16_mAd724_1 CB@16_mAd724_2 CB@16_mAd725_1 CB@16_mAd725_2 CB@16_mAd726_1 CB@16_mAd726_2 CB@16_mAd727_1 CB@16_mAd727_2 CB@16_mAd730_1 CB@16_mAd730_2 CB@16_mAd731_1 CB@16_mAd731_2 CB@16_mAd732_1 CB@16_mAd732_2 CB@16_mAd733_1 CB@16_mAd733_2 CB@16_mAd734_1 CB@16_mAd734_2 CB@16_mAd735_1 CB@16_mAd735_2 CB@16_mAd736_1 
+CB@16_mAd736_2 CB@16_mAd737_1 CB@16_mAd737_2 CB@16_mAd740_1 CB@16_mAd740_2 CB@16_mAd741_1 CB@16_mAd741_2 CB@16_mAd742_1 CB@16_mAd742_2 CB@16_mAd743_1 CB@16_mAd743_2 CB@16_mAd744_1 CB@16_mAd744_2 CB@16_mAd745_1 CB@16_mAd745_2 CB@16_mAd746_1 CB@16_mAd746_2 CB@16_mAd747_1 CB@16_mAd747_2 CB@16_mAd750_1 CB@16_mAd750_2 CB@16_mAd751_1 CB@16_mAd751_2 CB@16_mAd752_1 CB@16_mAd752_2 CB@16_mAd753_1 CB@16_mAd753_2 CB@16_mAd754_1 CB@16_mAd754_2 CB@16_mAd755_1 CB@16_mAd755_2 CB@16_mAd756_1 CB@16_mAd756_2 CB@16_mAd757_1 
+CB@16_mAd757_2 CB@16_mAd760_1 CB@16_mAd760_2 CB@16_mAd761_1 CB@16_mAd761_2 CB@16_mAd762_1 CB@16_mAd762_2 CB@16_mAd763_1 CB@16_mAd763_2 CB@16_mAd764_1 CB@16_mAd764_2 CB@16_mAd765_1 CB@16_mAd765_2 CB@16_mAd766_1 CB@16_mAd766_2 CB@16_mAd767_1 CB@16_mAd767_2 CB@16_mAd771_1 CB@16_mAd771_2 CB@16_mAd772_1 CB@16_mAd772_2 CB@16_mAd773_1 CB@16_mAd773_2 CB@16_mAd774_1 CB@16_mAd774_2 CB@16_mAd775_1 CB@16_mAd775_2 CB@16_mAd776_1 CB@16_mAd776_2 CB@16_mAd777_1 CB@16_mAd777_2 CB@16_X0 CB@16_X1 CB@16_X10 CB@16_X11 
+CB@16_X12 CB@16_X13 CB@16_X2 CB@16_X3 CB@16_X4 CB@16_X5 CB@16_X6 CB@16_X7 CB@16_X8 CB@16_X9 CB@16_Y1 CB@16_Y10 CB@16_Y11 CB@16_Y12 CB@16_Y2 CB@16_Y3 CB@16_Y4 CB@16_Y5 CB@16_Y6 CB@16_Y7 CB@16_Y8 CB@16_Y9 CB@16_Z1 CB@16_Z10 CB@16_Z11 CB@16_Z12 CB@16_Z2 CB@16_Z3 CB@16_Z4 CB@16_Z5 CB@16_Z6 CB@16_Z7 CB@16_Z8 CB@16_Z9 _5400TP094__CB
XCB@17 CB@17_K0 CB@17_K1 CB@17_K10 CB@17_K11 CB@17_K12 CB@17_K13 CB@17_K2 CB@17_K3 CB@17_K4 CB@17_K5 CB@17_K6 CB@17_K7 CB@17_K8 CB@17_K9 CB@17_mAd000_1 CB@17_mAd000_2 CB@17_mAd001_1 CB@17_mAd001_2 CB@17_mAd002_1 CB@17_mAd002_2 CB@17_mAd003_1 CB@17_mAd003_2 CB@17_mAd004_1 CB@17_mAd004_2 CB@17_mAd005_1 CB@17_mAd005_2 CB@17_mAd006_1 CB@17_mAd006_2 CB@17_mAd007_1 CB@17_mAd007_2 CB@17_mAd010_1 CB@17_mAd010_2 CB@17_mAd011_1 CB@17_mAd011_2 CB@17_mAd012_1 CB@17_mAd012_2 CB@17_mAd013_1 CB@17_mAd013_2 CB@17_mAd014_1 
+CB@17_mAd014_2 CB@17_mAd015_1 CB@17_mAd015_2 CB@17_mAd016_1 CB@17_mAd016_2 CB@17_mAd017_1 CB@17_mAd017_2 CB@17_mAd020_1 CB@17_mAd020_2 CB@17_mAd021_1 CB@17_mAd021_2 CB@17_mAd022_1 CB@17_mAd022_2 CB@17_mAd023_1 CB@17_mAd023_2 CB@17_mAd024_1 CB@17_mAd024_2 CB@17_mAd025_1 CB@17_mAd025_2 CB@17_mAd026_1 CB@17_mAd026_2 CB@17_mAd027_1 CB@17_mAd027_2 CB@17_mAd030_1 CB@17_mAd030_2 CB@17_mAd031_1 CB@17_mAd031_2 CB@17_mAd032_1 CB@17_mAd032_2 CB@17_mAd033_1 CB@17_mAd033_2 CB@17_mAd034_1 CB@17_mAd034_2 CB@17_mAd035_1 
+CB@17_mAd035_2 CB@17_mAd036_1 CB@17_mAd036_2 CB@17_mAd037_1 CB@17_mAd037_2 CB@17_mAd040_1 CB@17_mAd040_2 CB@17_mAd041_1 CB@17_mAd041_2 CB@17_mAd042_1 CB@17_mAd042_2 CB@17_mAd043_1 CB@17_mAd043_2 CB@17_mAd044_1 CB@17_mAd044_2 CB@17_mAd045_1 CB@17_mAd045_2 CB@17_mAd046_1 CB@17_mAd046_2 CB@17_mAd047_1 CB@17_mAd047_2 CB@17_mAd050_1 CB@17_mAd050_2 CB@17_mAd051_1 CB@17_mAd051_2 CB@17_mAd052_1 CB@17_mAd052_2 CB@17_mAd053_1 CB@17_mAd053_2 CB@17_mAd054_1 CB@17_mAd054_2 CB@17_mAd055_1 CB@17_mAd055_2 CB@17_mAd056_1 
+CB@17_mAd056_2 CB@17_mAd057_1 CB@17_mAd057_2 CB@17_mAd060_1 CB@17_mAd060_2 CB@17_mAd066_1 CB@17_mAd066_2 CB@17_mAd067_1 CB@17_mAd067_2 CB@17_mAd100_1 CB@17_mAd100_2 CB@17_mAd101_1 CB@17_mAd101_2 CB@17_mAd102_1 CB@17_mAd102_2 CB@17_mAd110_1 CB@17_mAd110_2 CB@17_mAd111_1 CB@17_mAd111_2 CB@17_mAd112_1 CB@17_mAd112_2 CB@17_mAd113_1 CB@17_mAd113_2 CB@17_mAd114_1 CB@17_mAd114_2 CB@17_mAd115_1 CB@17_mAd115_2 CB@17_mAd116_1 CB@17_mAd116_2 CB@17_mAd117_1 CB@17_mAd117_2 CB@17_mAd120_1 CB@17_mAd120_2 CB@17_mAd121_1 
+CB@17_mAd121_2 CB@17_mAd122_1 CB@17_mAd122_2 CB@17_mAd123_1 CB@17_mAd123_2 CB@17_mAd124_1 CB@17_mAd124_2 CB@17_mAd125_1 CB@17_mAd125_2 CB@17_mAd126_1 CB@17_mAd126_2 CB@17_mAd127_1 CB@17_mAd127_2 CB@17_mAd130_1 CB@17_mAd130_2 CB@17_mAd131_1 CB@17_mAd131_2 CB@17_mAd132_1 CB@17_mAd132_2 CB@17_mAd133_1 CB@17_mAd133_2 CB@17_mAd134_1 CB@17_mAd134_2 CB@17_mAd135_1 CB@17_mAd135_2 CB@17_mAd136_1 CB@17_mAd136_2 CB@17_mAd137_1 CB@17_mAd137_2 CB@17_mAd140_1 CB@17_mAd140_2 CB@17_mAd141_1 CB@17_mAd141_2 CB@17_mAd142_1 
+CB@17_mAd142_2 CB@17_mAd143_1 CB@17_mAd143_2 CB@17_mAd144_1 CB@17_mAd144_2 CB@17_mAd145_1 CB@17_mAd145_2 CB@17_mAd146_1 CB@17_mAd146_2 CB@17_mAd147_1 CB@17_mAd147_2 CB@17_mAd150_1 CB@17_mAd150_2 CB@17_mAd151_1 CB@17_mAd151_2 CB@17_mAd152_1 CB@17_mAd152_2 CB@17_mAd153_1 CB@17_mAd153_2 CB@17_mAd154_1 CB@17_mAd154_2 CB@17_mAd155_1 CB@17_mAd155_2 CB@17_mAd156_1 CB@17_mAd156_2 CB@17_mAd157_1 CB@17_mAd157_2 CB@17_mAd160_1 CB@17_mAd160_2 CB@17_mAd161_1 CB@17_mAd161_2 CB@17_mAd162_1 CB@17_mAd162_2 CB@17_mAd163_1 
+CB@17_mAd163_2 CB@17_mAd164_1 CB@17_mAd164_2 CB@17_mAd165_1 CB@17_mAd165_2 CB@17_mAd166_1 CB@17_mAd166_2 CB@17_mAd167_1 CB@17_mAd167_2 CB@17_mAd170_1 CB@17_mAd170_2 CB@17_mAd171_1 CB@17_mAd171_2 CB@17_mAd172_1 CB@17_mAd172_2 CB@17_mAd173_1 CB@17_mAd173_2 CB@17_mAd175_1 CB@17_mAd175_2 CB@17_mAd176_1 CB@17_mAd176_2 CB@17_mAd177_1 CB@17_mAd177_2 CB@17_mAd200_1 CB@17_mAd200_2 CB@17_mAd201_1 CB@17_mAd201_2 CB@17_mAd202_1 CB@17_mAd202_2 CB@17_mAd204_1 CB@17_mAd204_2 CB@17_mAd205_1 CB@17_mAd205_2 CB@17_mAd206_1 
+CB@17_mAd206_2 CB@17_mAd207_1 CB@17_mAd207_2 CB@17_mAd210_1 CB@17_mAd210_2 CB@17_mAd211_1 CB@17_mAd211_2 CB@17_mAd212_1 CB@17_mAd212_2 CB@17_mAd213_1 CB@17_mAd213_2 CB@17_mAd214_1 CB@17_mAd214_2 CB@17_mAd215_1 CB@17_mAd215_2 CB@17_mAd216_1 CB@17_mAd216_2 CB@17_mAd217_1 CB@17_mAd217_2 CB@17_mAd220_1 CB@17_mAd220_2 CB@17_mAd221_1 CB@17_mAd221_2 CB@17_mAd222_1 CB@17_mAd222_2 CB@17_mAd223_1 CB@17_mAd223_2 CB@17_mAd224_1 CB@17_mAd224_2 CB@17_mAd225_1 CB@17_mAd225_2 CB@17_mAd226_1 CB@17_mAd226_2 CB@17_mAd227_1 
+CB@17_mAd227_2 CB@17_mAd230_1 CB@17_mAd230_2 CB@17_mAd231_1 CB@17_mAd231_2 CB@17_mAd232_1 CB@17_mAd232_2 CB@17_mAd233_1 CB@17_mAd233_2 CB@17_mAd234_1 CB@17_mAd234_2 CB@17_mAd235_1 CB@17_mAd235_2 CB@17_mAd236_1 CB@17_mAd236_2 CB@17_mAd237_1 CB@17_mAd237_2 CB@17_mAd240_1 CB@17_mAd240_2 CB@17_mAd241_1 CB@17_mAd241_2 CB@17_mAd242_1 CB@17_mAd242_2 CB@17_mAd243_1 CB@17_mAd243_2 CB@17_mAd244_1 CB@17_mAd244_2 CB@17_mAd245_1 CB@17_mAd245_2 CB@17_mAd246_1 CB@17_mAd246_2 CB@17_mAd247_1 CB@17_mAd247_2 CB@17_mAd250_1 
+CB@17_mAd250_2 CB@17_mAd251_1 CB@17_mAd251_2 CB@17_mAd252_1 CB@17_mAd252_2 CB@17_mAd253_1 CB@17_mAd253_2 CB@17_mAd254_1 CB@17_mAd254_2 CB@17_mAd255_1 CB@17_mAd255_2 CB@17_mAd256_1 CB@17_mAd256_2 CB@17_mAd257_1 CB@17_mAd257_2 CB@17_mAd260_1 CB@17_mAd260_2 CB@17_mAd261_1 CB@17_mAd261_2 CB@17_mAd262_1 CB@17_mAd262_2 CB@17_mAd263_1 CB@17_mAd263_2 CB@17_mAd264_1 CB@17_mAd264_2 CB@17_mAd265_1 CB@17_mAd265_2 CB@17_mAd266_1 CB@17_mAd266_2 CB@17_mAd267_1 CB@17_mAd267_2 CB@17_mAd275_1 CB@17_mAd275_2 CB@17_mAd276_1 
+CB@17_mAd276_2 CB@17_mAd277_1 CB@17_mAd277_2 CB@17_mAd300_1 CB@17_mAd300_2 CB@17_mAd310_1 CB@17_mAd310_2 CB@17_mAd311_1 CB@17_mAd311_2 CB@17_mAd317_1 CB@17_mAd317_2 CB@17_mAd320_1 CB@17_mAd320_2 CB@17_mAd321_1 CB@17_mAd321_2 CB@17_mAd322_1 CB@17_mAd322_2 CB@17_mAd323_1 CB@17_mAd323_2 CB@17_mAd324_1 CB@17_mAd324_2 CB@17_mAd325_1 CB@17_mAd325_2 CB@17_mAd326_1 CB@17_mAd326_2 CB@17_mAd327_1 CB@17_mAd327_2 CB@17_mAd330_1 CB@17_mAd330_2 CB@17_mAd331_1 CB@17_mAd331_2 CB@17_mAd332_1 CB@17_mAd332_2 CB@17_mAd333_1 
+CB@17_mAd333_2 CB@17_mAd334_1 CB@17_mAd334_2 CB@17_mAd335_1 CB@17_mAd335_2 CB@17_mAd336_1 CB@17_mAd336_2 CB@17_mAd337_1 CB@17_mAd337_2 CB@17_mAd340_1 CB@17_mAd340_2 CB@17_mAd341_1 CB@17_mAd341_2 CB@17_mAd342_1 CB@17_mAd342_2 CB@17_mAd343_1 CB@17_mAd343_2 CB@17_mAd344_1 CB@17_mAd344_2 CB@17_mAd345_1 CB@17_mAd345_2 CB@17_mAd346_1 CB@17_mAd346_2 CB@17_mAd347_1 CB@17_mAd347_2 CB@17_mAd350_1 CB@17_mAd350_2 CB@17_mAd351_1 CB@17_mAd351_2 CB@17_mAd352_1 CB@17_mAd352_2 CB@17_mAd353_1 CB@17_mAd353_2 CB@17_mAd354_1 
+CB@17_mAd354_2 CB@17_mAd355_1 CB@17_mAd355_2 CB@17_mAd356_1 CB@17_mAd356_2 CB@17_mAd357_1 CB@17_mAd357_2 CB@17_mAd360_1 CB@17_mAd360_2 CB@17_mAd361_1 CB@17_mAd361_2 CB@17_mAd362_1 CB@17_mAd362_2 CB@17_mAd363_1 CB@17_mAd363_2 CB@17_mAd364_1 CB@17_mAd364_2 CB@17_mAd365_1 CB@17_mAd365_2 CB@17_mAd366_1 CB@17_mAd366_2 CB@17_mAd367_1 CB@17_mAd367_2 CB@17_mAd371_1 CB@17_mAd371_2 CB@17_mAd372_1 CB@17_mAd372_2 CB@17_mAd373_1 CB@17_mAd373_2 CB@17_mAd374_1 CB@17_mAd374_2 CB@17_mAd375_1 CB@17_mAd375_2 CB@17_mAd376_1 
+CB@17_mAd376_2 CB@17_mAd377_1 CB@17_mAd377_2 CB@17_mAd400_1 CB@17_mAd400_2 CB@17_mAd401_1 CB@17_mAd401_2 CB@17_mAd402_1 CB@17_mAd402_2 CB@17_mAd403_1 CB@17_mAd403_2 CB@17_mAd404_1 CB@17_mAd404_2 CB@17_mAd405_1 CB@17_mAd405_2 CB@17_mAd406_1 CB@17_mAd406_2 CB@17_mAd407_1 CB@17_mAd407_2 CB@17_mAd410_1 CB@17_mAd410_2 CB@17_mAd411_1 CB@17_mAd411_2 CB@17_mAd412_1 CB@17_mAd412_2 CB@17_mAd413_1 CB@17_mAd413_2 CB@17_mAd414_1 CB@17_mAd414_2 CB@17_mAd415_1 CB@17_mAd415_2 CB@17_mAd416_1 CB@17_mAd416_2 CB@17_mAd417_1 
+CB@17_mAd417_2 CB@17_mAd420_1 CB@17_mAd420_2 CB@17_mAd421_1 CB@17_mAd421_2 CB@17_mAd422_1 CB@17_mAd422_2 CB@17_mAd423_1 CB@17_mAd423_2 CB@17_mAd424_1 CB@17_mAd424_2 CB@17_mAd425_1 CB@17_mAd425_2 CB@17_mAd426_1 CB@17_mAd426_2 CB@17_mAd427_1 CB@17_mAd427_2 CB@17_mAd430_1 CB@17_mAd430_2 CB@17_mAd431_1 CB@17_mAd431_2 CB@17_mAd432_1 CB@17_mAd432_2 CB@17_mAd433_1 CB@17_mAd433_2 CB@17_mAd434_1 CB@17_mAd434_2 CB@17_mAd435_1 CB@17_mAd435_2 CB@17_mAd436_1 CB@17_mAd436_2 CB@17_mAd437_1 CB@17_mAd437_2 CB@17_mAd440_1 
+CB@17_mAd440_2 CB@17_mAd441_1 CB@17_mAd441_2 CB@17_mAd442_1 CB@17_mAd442_2 CB@17_mAd443_1 CB@17_mAd443_2 CB@17_mAd444_1 CB@17_mAd444_2 CB@17_mAd445_1 CB@17_mAd445_2 CB@17_mAd446_1 CB@17_mAd446_2 CB@17_mAd447_1 CB@17_mAd447_2 CB@17_mAd450_1 CB@17_mAd450_2 CB@17_mAd451_1 CB@17_mAd451_2 CB@17_mAd452_1 CB@17_mAd452_2 CB@17_mAd453_1 CB@17_mAd453_2 CB@17_mAd454_1 CB@17_mAd454_2 CB@17_mAd455_1 CB@17_mAd455_2 CB@17_mAd456_1 CB@17_mAd456_2 CB@17_mAd457_1 CB@17_mAd457_2 CB@17_mAd460_1 CB@17_mAd460_2 CB@17_mAd466_1 
+CB@17_mAd466_2 CB@17_mAd467_1 CB@17_mAd467_2 CB@17_mAd500_1 CB@17_mAd500_2 CB@17_mAd501_1 CB@17_mAd501_2 CB@17_mAd502_1 CB@17_mAd502_2 CB@17_mAd508_1 CB@17_mAd508_2 CB@17_mAd509_1 CB@17_mAd509_2 CB@17_mAd512_1 CB@17_mAd512_2 CB@17_mAd513_1 CB@17_mAd513_2 CB@17_mAd514_1 CB@17_mAd514_2 CB@17_mAd515_1 CB@17_mAd515_2 CB@17_mAd516_1 CB@17_mAd516_2 CB@17_mAd517_1 CB@17_mAd517_2 CB@17_mAd520_1 CB@17_mAd520_2 CB@17_mAd521_1 CB@17_mAd521_2 CB@17_mAd522_1 CB@17_mAd522_2 CB@17_mAd523_1 CB@17_mAd523_2 CB@17_mAd524_1 
+CB@17_mAd524_2 CB@17_mAd525_1 CB@17_mAd525_2 CB@17_mAd526_1 CB@17_mAd526_2 CB@17_mAd527_1 CB@17_mAd527_2 CB@17_mAd530_1 CB@17_mAd530_2 CB@17_mAd531_1 CB@17_mAd531_2 CB@17_mAd532_1 CB@17_mAd532_2 CB@17_mAd533_1 CB@17_mAd533_2 CB@17_mAd534_1 CB@17_mAd534_2 CB@17_mAd535_1 CB@17_mAd535_2 CB@17_mAd536_1 CB@17_mAd536_2 CB@17_mAd537_1 CB@17_mAd537_2 CB@17_mAd540_1 CB@17_mAd540_2 CB@17_mAd541_1 CB@17_mAd541_2 CB@17_mAd542_1 CB@17_mAd542_2 CB@17_mAd543_1 CB@17_mAd543_2 CB@17_mAd544_1 CB@17_mAd544_2 CB@17_mAd545_1 
+CB@17_mAd545_2 CB@17_mAd546_1 CB@17_mAd546_2 CB@17_mAd547_1 CB@17_mAd547_2 CB@17_mAd550_1 CB@17_mAd550_2 CB@17_mAd551_1 CB@17_mAd551_2 CB@17_mAd552_1 CB@17_mAd552_2 CB@17_mAd553_1 CB@17_mAd553_2 CB@17_mAd554_1 CB@17_mAd554_2 CB@17_mAd555_1 CB@17_mAd555_2 CB@17_mAd556_1 CB@17_mAd556_2 CB@17_mAd557_1 CB@17_mAd557_2 CB@17_mAd560_1 CB@17_mAd560_2 CB@17_mAd561_1 CB@17_mAd561_2 CB@17_mAd562_1 CB@17_mAd562_2 CB@17_mAd563_1 CB@17_mAd563_2 CB@17_mAd564_1 CB@17_mAd564_2 CB@17_mAd565_1 CB@17_mAd565_2 CB@17_mAd566_1 
+CB@17_mAd566_2 CB@17_mAd567_1 CB@17_mAd567_2 CB@17_mAd570_1 CB@17_mAd570_2 CB@17_mAd571_1 CB@17_mAd571_2 CB@17_mAd572_1 CB@17_mAd572_2 CB@17_mAd573_1 CB@17_mAd573_2 CB@17_mAd575_1 CB@17_mAd575_2 CB@17_mAd576_1 CB@17_mAd576_2 CB@17_mAd577_1 CB@17_mAd577_2 CB@17_mAd600_1 CB@17_mAd600_2 CB@17_mAd601_1 CB@17_mAd601_2 CB@17_mAd602_1 CB@17_mAd602_2 CB@17_mAd604_1 CB@17_mAd604_2 CB@17_mAd605_1 CB@17_mAd605_2 CB@17_mAd606_1 CB@17_mAd606_2 CB@17_mAd607_1 CB@17_mAd607_2 CB@17_mAd610_1 CB@17_mAd610_2 CB@17_mAd611_1 
+CB@17_mAd611_2 CB@17_mAd612_1 CB@17_mAd612_2 CB@17_mAd613_1 CB@17_mAd613_2 CB@17_mAd614_1 CB@17_mAd614_2 CB@17_mAd615_1 CB@17_mAd615_2 CB@17_mAd616_1 CB@17_mAd616_2 CB@17_mAd617_1 CB@17_mAd617_2 CB@17_mAd620_1 CB@17_mAd620_2 CB@17_mAd621_1 CB@17_mAd621_2 CB@17_mAd622_1 CB@17_mAd622_2 CB@17_mAd623_1 CB@17_mAd623_2 CB@17_mAd624_1 CB@17_mAd624_2 CB@17_mAd625_1 CB@17_mAd625_2 CB@17_mAd626_1 CB@17_mAd626_2 CB@17_mAd627_1 CB@17_mAd627_2 CB@17_mAd630_1 CB@17_mAd630_2 CB@17_mAd631_1 CB@17_mAd631_2 CB@17_mAd632_1 
+CB@17_mAd632_2 CB@17_mAd633_1 CB@17_mAd633_2 CB@17_mAd634_1 CB@17_mAd634_2 CB@17_mAd635_1 CB@17_mAd635_2 CB@17_mAd636_1 CB@17_mAd636_2 CB@17_mAd637_1 CB@17_mAd637_2 CB@17_mAd640_1 CB@17_mAd640_2 CB@17_mAd641_1 CB@17_mAd641_2 CB@17_mAd642_1 CB@17_mAd642_2 CB@17_mAd643_1 CB@17_mAd643_2 CB@17_mAd644_1 CB@17_mAd644_2 CB@17_mAd645_1 CB@17_mAd645_2 CB@17_mAd646_1 CB@17_mAd646_2 CB@17_mAd647_1 CB@17_mAd647_2 CB@17_mAd650_1 CB@17_mAd650_2 CB@17_mAd651_1 CB@17_mAd651_2 CB@17_mAd652_1 CB@17_mAd652_2 CB@17_mAd653_1 
+CB@17_mAd653_2 CB@17_mAd654_1 CB@17_mAd654_2 CB@17_mAd655_1 CB@17_mAd655_2 CB@17_mAd656_1 CB@17_mAd656_2 CB@17_mAd657_1 CB@17_mAd657_2 CB@17_mAd660_1 CB@17_mAd660_2 CB@17_mAd661_1 CB@17_mAd661_2 CB@17_mAd662_1 CB@17_mAd662_2 CB@17_mAd663_1 CB@17_mAd663_2 CB@17_mAd664_1 CB@17_mAd664_2 CB@17_mAd665_1 CB@17_mAd665_2 CB@17_mAd666_1 CB@17_mAd666_2 CB@17_mAd667_1 CB@17_mAd667_2 CB@17_mAd675_1 CB@17_mAd675_2 CB@17_mAd676_1 CB@17_mAd676_2 CB@17_mAd677_1 CB@17_mAd677_2 CB@17_mAd700_1 CB@17_mAd700_2 CB@17_mAd710_1 
+CB@17_mAd710_2 CB@17_mAd711_1 CB@17_mAd711_2 CB@17_mAd717_1 CB@17_mAd717_2 CB@17_mAd720_1 CB@17_mAd720_2 CB@17_mAd721_1 CB@17_mAd721_2 CB@17_mAd722_1 CB@17_mAd722_2 CB@17_mAd723_1 CB@17_mAd723_2 CB@17_mAd724_1 CB@17_mAd724_2 CB@17_mAd725_1 CB@17_mAd725_2 CB@17_mAd726_1 CB@17_mAd726_2 CB@17_mAd727_1 CB@17_mAd727_2 CB@17_mAd730_1 CB@17_mAd730_2 CB@17_mAd731_1 CB@17_mAd731_2 CB@17_mAd732_1 CB@17_mAd732_2 CB@17_mAd733_1 CB@17_mAd733_2 CB@17_mAd734_1 CB@17_mAd734_2 CB@17_mAd735_1 CB@17_mAd735_2 CB@17_mAd736_1 
+CB@17_mAd736_2 CB@17_mAd737_1 CB@17_mAd737_2 CB@17_mAd740_1 CB@17_mAd740_2 CB@17_mAd741_1 CB@17_mAd741_2 CB@17_mAd742_1 CB@17_mAd742_2 CB@17_mAd743_1 CB@17_mAd743_2 CB@17_mAd744_1 CB@17_mAd744_2 CB@17_mAd745_1 CB@17_mAd745_2 CB@17_mAd746_1 CB@17_mAd746_2 CB@17_mAd747_1 CB@17_mAd747_2 CB@17_mAd750_1 CB@17_mAd750_2 CB@17_mAd751_1 CB@17_mAd751_2 CB@17_mAd752_1 CB@17_mAd752_2 CB@17_mAd753_1 CB@17_mAd753_2 CB@17_mAd754_1 CB@17_mAd754_2 CB@17_mAd755_1 CB@17_mAd755_2 CB@17_mAd756_1 CB@17_mAd756_2 CB@17_mAd757_1 
+CB@17_mAd757_2 CB@17_mAd760_1 CB@17_mAd760_2 CB@17_mAd761_1 CB@17_mAd761_2 CB@17_mAd762_1 CB@17_mAd762_2 CB@17_mAd763_1 CB@17_mAd763_2 CB@17_mAd764_1 CB@17_mAd764_2 CB@17_mAd765_1 CB@17_mAd765_2 CB@17_mAd766_1 CB@17_mAd766_2 CB@17_mAd767_1 CB@17_mAd767_2 CB@17_mAd771_1 CB@17_mAd771_2 CB@17_mAd772_1 CB@17_mAd772_2 CB@17_mAd773_1 CB@17_mAd773_2 CB@17_mAd774_1 CB@17_mAd774_2 CB@17_mAd775_1 CB@17_mAd775_2 CB@17_mAd776_1 CB@17_mAd776_2 CB@17_mAd777_1 CB@17_mAd777_2 CB@17_X0 CB@17_X1 CB@17_X10 CB@17_X11 
+CB@17_X12 CB@17_X13 CB@17_X2 CB@17_X3 CB@17_X4 CB@17_X5 CB@17_X6 CB@17_X7 CB@17_X8 CB@17_X9 CB@17_Y1 CB@17_Y10 CB@17_Y11 CB@17_Y12 CB@17_Y2 CB@17_Y3 CB@17_Y4 CB@17_Y5 CB@17_Y6 CB@17_Y7 CB@17_Y8 CB@17_Y9 CB@17_Z1 CB@17_Z10 CB@17_Z11 CB@17_Z12 CB@17_Z2 CB@17_Z3 CB@17_Z4 CB@17_Z5 CB@17_Z6 CB@17_Z7 CB@17_Z8 CB@17_Z9 _5400TP094__CB
XCB@18 CB@18_K0 CB@18_K1 CB@18_K10 CB@18_K11 CB@18_K12 CB@18_K13 CB@18_K2 CB@18_K3 CB@18_K4 CB@18_K5 CB@18_K6 CB@18_K7 CB@18_K8 CB@18_K9 CB@18_mAd000_1 CB@18_mAd000_2 CB@18_mAd001_1 CB@18_mAd001_2 CB@18_mAd002_1 CB@18_mAd002_2 CB@18_mAd003_1 CB@18_mAd003_2 CB@18_mAd004_1 CB@18_mAd004_2 CB@18_mAd005_1 CB@18_mAd005_2 CB@18_mAd006_1 CB@18_mAd006_2 CB@18_mAd007_1 CB@18_mAd007_2 CB@18_mAd010_1 CB@18_mAd010_2 CB@18_mAd011_1 CB@18_mAd011_2 CB@18_mAd012_1 CB@18_mAd012_2 CB@18_mAd013_1 CB@18_mAd013_2 CB@18_mAd014_1 
+CB@18_mAd014_2 CB@18_mAd015_1 CB@18_mAd015_2 CB@18_mAd016_1 CB@18_mAd016_2 CB@18_mAd017_1 CB@18_mAd017_2 CB@18_mAd020_1 CB@18_mAd020_2 CB@18_mAd021_1 CB@18_mAd021_2 CB@18_mAd022_1 CB@18_mAd022_2 CB@18_mAd023_1 CB@18_mAd023_2 CB@18_mAd024_1 CB@18_mAd024_2 CB@18_mAd025_1 CB@18_mAd025_2 CB@18_mAd026_1 CB@18_mAd026_2 CB@18_mAd027_1 CB@18_mAd027_2 CB@18_mAd030_1 CB@18_mAd030_2 CB@18_mAd031_1 CB@18_mAd031_2 CB@18_mAd032_1 CB@18_mAd032_2 CB@18_mAd033_1 CB@18_mAd033_2 CB@18_mAd034_1 CB@18_mAd034_2 CB@18_mAd035_1 
+CB@18_mAd035_2 CB@18_mAd036_1 CB@18_mAd036_2 CB@18_mAd037_1 CB@18_mAd037_2 CB@18_mAd040_1 CB@18_mAd040_2 CB@18_mAd041_1 CB@18_mAd041_2 CB@18_mAd042_1 CB@18_mAd042_2 CB@18_mAd043_1 CB@18_mAd043_2 CB@18_mAd044_1 CB@18_mAd044_2 CB@18_mAd045_1 CB@18_mAd045_2 CB@18_mAd046_1 CB@18_mAd046_2 CB@18_mAd047_1 CB@18_mAd047_2 CB@18_mAd050_1 CB@18_mAd050_2 CB@18_mAd051_1 CB@18_mAd051_2 CB@18_mAd052_1 CB@18_mAd052_2 CB@18_mAd053_1 CB@18_mAd053_2 CB@18_mAd054_1 CB@18_mAd054_2 CB@18_mAd055_1 CB@18_mAd055_2 CB@18_mAd056_1 
+CB@18_mAd056_2 CB@18_mAd057_1 CB@18_mAd057_2 CB@18_mAd060_1 CB@18_mAd060_2 CB@18_mAd066_1 CB@18_mAd066_2 CB@18_mAd067_1 CB@18_mAd067_2 CB@18_mAd100_1 CB@18_mAd100_2 CB@18_mAd101_1 CB@18_mAd101_2 CB@18_mAd102_1 CB@18_mAd102_2 CB@18_mAd110_1 CB@18_mAd110_2 CB@18_mAd111_1 CB@18_mAd111_2 CB@18_mAd112_1 CB@18_mAd112_2 CB@18_mAd113_1 CB@18_mAd113_2 CB@18_mAd114_1 CB@18_mAd114_2 CB@18_mAd115_1 CB@18_mAd115_2 CB@18_mAd116_1 CB@18_mAd116_2 CB@18_mAd117_1 CB@18_mAd117_2 CB@18_mAd120_1 CB@18_mAd120_2 CB@18_mAd121_1 
+CB@18_mAd121_2 CB@18_mAd122_1 CB@18_mAd122_2 CB@18_mAd123_1 CB@18_mAd123_2 CB@18_mAd124_1 CB@18_mAd124_2 CB@18_mAd125_1 CB@18_mAd125_2 CB@18_mAd126_1 CB@18_mAd126_2 CB@18_mAd127_1 CB@18_mAd127_2 CB@18_mAd130_1 CB@18_mAd130_2 CB@18_mAd131_1 CB@18_mAd131_2 CB@18_mAd132_1 CB@18_mAd132_2 CB@18_mAd133_1 CB@18_mAd133_2 CB@18_mAd134_1 CB@18_mAd134_2 CB@18_mAd135_1 CB@18_mAd135_2 CB@18_mAd136_1 CB@18_mAd136_2 CB@18_mAd137_1 CB@18_mAd137_2 CB@18_mAd140_1 CB@18_mAd140_2 CB@18_mAd141_1 CB@18_mAd141_2 CB@18_mAd142_1 
+CB@18_mAd142_2 CB@18_mAd143_1 CB@18_mAd143_2 CB@18_mAd144_1 CB@18_mAd144_2 CB@18_mAd145_1 CB@18_mAd145_2 CB@18_mAd146_1 CB@18_mAd146_2 CB@18_mAd147_1 CB@18_mAd147_2 CB@18_mAd150_1 CB@18_mAd150_2 CB@18_mAd151_1 CB@18_mAd151_2 CB@18_mAd152_1 CB@18_mAd152_2 CB@18_mAd153_1 CB@18_mAd153_2 CB@18_mAd154_1 CB@18_mAd154_2 CB@18_mAd155_1 CB@18_mAd155_2 CB@18_mAd156_1 CB@18_mAd156_2 CB@18_mAd157_1 CB@18_mAd157_2 CB@18_mAd160_1 CB@18_mAd160_2 CB@18_mAd161_1 CB@18_mAd161_2 CB@18_mAd162_1 CB@18_mAd162_2 CB@18_mAd163_1 
+CB@18_mAd163_2 CB@18_mAd164_1 CB@18_mAd164_2 CB@18_mAd165_1 CB@18_mAd165_2 CB@18_mAd166_1 CB@18_mAd166_2 CB@18_mAd167_1 CB@18_mAd167_2 CB@18_mAd170_1 CB@18_mAd170_2 CB@18_mAd171_1 CB@18_mAd171_2 CB@18_mAd172_1 CB@18_mAd172_2 CB@18_mAd173_1 CB@18_mAd173_2 CB@18_mAd175_1 CB@18_mAd175_2 CB@18_mAd176_1 CB@18_mAd176_2 CB@18_mAd177_1 CB@18_mAd177_2 CB@18_mAd200_1 CB@18_mAd200_2 CB@18_mAd201_1 CB@18_mAd201_2 CB@18_mAd202_1 CB@18_mAd202_2 CB@18_mAd204_1 CB@18_mAd204_2 CB@18_mAd205_1 CB@18_mAd205_2 CB@18_mAd206_1 
+CB@18_mAd206_2 CB@18_mAd207_1 CB@18_mAd207_2 CB@18_mAd210_1 CB@18_mAd210_2 CB@18_mAd211_1 CB@18_mAd211_2 CB@18_mAd212_1 CB@18_mAd212_2 CB@18_mAd213_1 CB@18_mAd213_2 CB@18_mAd214_1 CB@18_mAd214_2 CB@18_mAd215_1 CB@18_mAd215_2 CB@18_mAd216_1 CB@18_mAd216_2 CB@18_mAd217_1 CB@18_mAd217_2 CB@18_mAd220_1 CB@18_mAd220_2 CB@18_mAd221_1 CB@18_mAd221_2 CB@18_mAd222_1 CB@18_mAd222_2 CB@18_mAd223_1 CB@18_mAd223_2 CB@18_mAd224_1 CB@18_mAd224_2 CB@18_mAd225_1 CB@18_mAd225_2 CB@18_mAd226_1 CB@18_mAd226_2 CB@18_mAd227_1 
+CB@18_mAd227_2 CB@18_mAd230_1 CB@18_mAd230_2 CB@18_mAd231_1 CB@18_mAd231_2 CB@18_mAd232_1 CB@18_mAd232_2 CB@18_mAd233_1 CB@18_mAd233_2 CB@18_mAd234_1 CB@18_mAd234_2 CB@18_mAd235_1 CB@18_mAd235_2 CB@18_mAd236_1 CB@18_mAd236_2 CB@18_mAd237_1 CB@18_mAd237_2 CB@18_mAd240_1 CB@18_mAd240_2 CB@18_mAd241_1 CB@18_mAd241_2 CB@18_mAd242_1 CB@18_mAd242_2 CB@18_mAd243_1 CB@18_mAd243_2 CB@18_mAd244_1 CB@18_mAd244_2 CB@18_mAd245_1 CB@18_mAd245_2 CB@18_mAd246_1 CB@18_mAd246_2 CB@18_mAd247_1 CB@18_mAd247_2 CB@18_mAd250_1 
+CB@18_mAd250_2 CB@18_mAd251_1 CB@18_mAd251_2 CB@18_mAd252_1 CB@18_mAd252_2 CB@18_mAd253_1 CB@18_mAd253_2 CB@18_mAd254_1 CB@18_mAd254_2 CB@18_mAd255_1 CB@18_mAd255_2 CB@18_mAd256_1 CB@18_mAd256_2 CB@18_mAd257_1 CB@18_mAd257_2 CB@18_mAd260_1 CB@18_mAd260_2 CB@18_mAd261_1 CB@18_mAd261_2 CB@18_mAd262_1 CB@18_mAd262_2 CB@18_mAd263_1 CB@18_mAd263_2 CB@18_mAd264_1 CB@18_mAd264_2 CB@18_mAd265_1 CB@18_mAd265_2 CB@18_mAd266_1 CB@18_mAd266_2 CB@18_mAd267_1 CB@18_mAd267_2 CB@18_mAd275_1 CB@18_mAd275_2 CB@18_mAd276_1 
+CB@18_mAd276_2 CB@18_mAd277_1 CB@18_mAd277_2 CB@18_mAd300_1 CB@18_mAd300_2 CB@18_mAd310_1 CB@18_mAd310_2 CB@18_mAd311_1 CB@18_mAd311_2 CB@18_mAd317_1 CB@18_mAd317_2 CB@18_mAd320_1 CB@18_mAd320_2 CB@18_mAd321_1 CB@18_mAd321_2 CB@18_mAd322_1 CB@18_mAd322_2 CB@18_mAd323_1 CB@18_mAd323_2 CB@18_mAd324_1 CB@18_mAd324_2 CB@18_mAd325_1 CB@18_mAd325_2 CB@18_mAd326_1 CB@18_mAd326_2 CB@18_mAd327_1 CB@18_mAd327_2 CB@18_mAd330_1 CB@18_mAd330_2 CB@18_mAd331_1 CB@18_mAd331_2 CB@18_mAd332_1 CB@18_mAd332_2 CB@18_mAd333_1 
+CB@18_mAd333_2 CB@18_mAd334_1 CB@18_mAd334_2 CB@18_mAd335_1 CB@18_mAd335_2 CB@18_mAd336_1 CB@18_mAd336_2 CB@18_mAd337_1 CB@18_mAd337_2 CB@18_mAd340_1 CB@18_mAd340_2 CB@18_mAd341_1 CB@18_mAd341_2 CB@18_mAd342_1 CB@18_mAd342_2 CB@18_mAd343_1 CB@18_mAd343_2 CB@18_mAd344_1 CB@18_mAd344_2 CB@18_mAd345_1 CB@18_mAd345_2 CB@18_mAd346_1 CB@18_mAd346_2 CB@18_mAd347_1 CB@18_mAd347_2 CB@18_mAd350_1 CB@18_mAd350_2 CB@18_mAd351_1 CB@18_mAd351_2 CB@18_mAd352_1 CB@18_mAd352_2 CB@18_mAd353_1 CB@18_mAd353_2 CB@18_mAd354_1 
+CB@18_mAd354_2 CB@18_mAd355_1 CB@18_mAd355_2 CB@18_mAd356_1 CB@18_mAd356_2 CB@18_mAd357_1 CB@18_mAd357_2 CB@18_mAd360_1 CB@18_mAd360_2 CB@18_mAd361_1 CB@18_mAd361_2 CB@18_mAd362_1 CB@18_mAd362_2 CB@18_mAd363_1 CB@18_mAd363_2 CB@18_mAd364_1 CB@18_mAd364_2 CB@18_mAd365_1 CB@18_mAd365_2 CB@18_mAd366_1 CB@18_mAd366_2 CB@18_mAd367_1 CB@18_mAd367_2 CB@18_mAd371_1 CB@18_mAd371_2 CB@18_mAd372_1 CB@18_mAd372_2 CB@18_mAd373_1 CB@18_mAd373_2 CB@18_mAd374_1 CB@18_mAd374_2 CB@18_mAd375_1 CB@18_mAd375_2 CB@18_mAd376_1 
+CB@18_mAd376_2 CB@18_mAd377_1 CB@18_mAd377_2 CB@18_mAd400_1 CB@18_mAd400_2 CB@18_mAd401_1 CB@18_mAd401_2 CB@18_mAd402_1 CB@18_mAd402_2 CB@18_mAd403_1 CB@18_mAd403_2 CB@18_mAd404_1 CB@18_mAd404_2 CB@18_mAd405_1 CB@18_mAd405_2 CB@18_mAd406_1 CB@18_mAd406_2 CB@18_mAd407_1 CB@18_mAd407_2 CB@18_mAd410_1 CB@18_mAd410_2 CB@18_mAd411_1 CB@18_mAd411_2 CB@18_mAd412_1 CB@18_mAd412_2 CB@18_mAd413_1 CB@18_mAd413_2 CB@18_mAd414_1 CB@18_mAd414_2 CB@18_mAd415_1 CB@18_mAd415_2 CB@18_mAd416_1 CB@18_mAd416_2 CB@18_mAd417_1 
+CB@18_mAd417_2 CB@18_mAd420_1 CB@18_mAd420_2 CB@18_mAd421_1 CB@18_mAd421_2 CB@18_mAd422_1 CB@18_mAd422_2 CB@18_mAd423_1 CB@18_mAd423_2 CB@18_mAd424_1 CB@18_mAd424_2 CB@18_mAd425_1 CB@18_mAd425_2 CB@18_mAd426_1 CB@18_mAd426_2 CB@18_mAd427_1 CB@18_mAd427_2 CB@18_mAd430_1 CB@18_mAd430_2 CB@18_mAd431_1 CB@18_mAd431_2 CB@18_mAd432_1 CB@18_mAd432_2 CB@18_mAd433_1 CB@18_mAd433_2 CB@18_mAd434_1 CB@18_mAd434_2 CB@18_mAd435_1 CB@18_mAd435_2 CB@18_mAd436_1 CB@18_mAd436_2 CB@18_mAd437_1 CB@18_mAd437_2 CB@18_mAd440_1 
+CB@18_mAd440_2 CB@18_mAd441_1 CB@18_mAd441_2 CB@18_mAd442_1 CB@18_mAd442_2 CB@18_mAd443_1 CB@18_mAd443_2 CB@18_mAd444_1 CB@18_mAd444_2 CB@18_mAd445_1 CB@18_mAd445_2 CB@18_mAd446_1 CB@18_mAd446_2 CB@18_mAd447_1 CB@18_mAd447_2 CB@18_mAd450_1 CB@18_mAd450_2 CB@18_mAd451_1 CB@18_mAd451_2 CB@18_mAd452_1 CB@18_mAd452_2 CB@18_mAd453_1 CB@18_mAd453_2 CB@18_mAd454_1 CB@18_mAd454_2 CB@18_mAd455_1 CB@18_mAd455_2 CB@18_mAd456_1 CB@18_mAd456_2 CB@18_mAd457_1 CB@18_mAd457_2 CB@18_mAd460_1 CB@18_mAd460_2 CB@18_mAd466_1 
+CB@18_mAd466_2 CB@18_mAd467_1 CB@18_mAd467_2 CB@18_mAd500_1 CB@18_mAd500_2 CB@18_mAd501_1 CB@18_mAd501_2 CB@18_mAd502_1 CB@18_mAd502_2 CB@18_mAd508_1 CB@18_mAd508_2 CB@18_mAd509_1 CB@18_mAd509_2 CB@18_mAd512_1 CB@18_mAd512_2 CB@18_mAd513_1 CB@18_mAd513_2 CB@18_mAd514_1 CB@18_mAd514_2 CB@18_mAd515_1 CB@18_mAd515_2 CB@18_mAd516_1 CB@18_mAd516_2 CB@18_mAd517_1 CB@18_mAd517_2 CB@18_mAd520_1 CB@18_mAd520_2 CB@18_mAd521_1 CB@18_mAd521_2 CB@18_mAd522_1 CB@18_mAd522_2 CB@18_mAd523_1 CB@18_mAd523_2 CB@18_mAd524_1 
+CB@18_mAd524_2 CB@18_mAd525_1 CB@18_mAd525_2 CB@18_mAd526_1 CB@18_mAd526_2 CB@18_mAd527_1 CB@18_mAd527_2 CB@18_mAd530_1 CB@18_mAd530_2 CB@18_mAd531_1 CB@18_mAd531_2 CB@18_mAd532_1 CB@18_mAd532_2 CB@18_mAd533_1 CB@18_mAd533_2 CB@18_mAd534_1 CB@18_mAd534_2 CB@18_mAd535_1 CB@18_mAd535_2 CB@18_mAd536_1 CB@18_mAd536_2 CB@18_mAd537_1 CB@18_mAd537_2 CB@18_mAd540_1 CB@18_mAd540_2 CB@18_mAd541_1 CB@18_mAd541_2 CB@18_mAd542_1 CB@18_mAd542_2 CB@18_mAd543_1 CB@18_mAd543_2 CB@18_mAd544_1 CB@18_mAd544_2 CB@18_mAd545_1 
+CB@18_mAd545_2 CB@18_mAd546_1 CB@18_mAd546_2 CB@18_mAd547_1 CB@18_mAd547_2 CB@18_mAd550_1 CB@18_mAd550_2 CB@18_mAd551_1 CB@18_mAd551_2 CB@18_mAd552_1 CB@18_mAd552_2 CB@18_mAd553_1 CB@18_mAd553_2 CB@18_mAd554_1 CB@18_mAd554_2 CB@18_mAd555_1 CB@18_mAd555_2 CB@18_mAd556_1 CB@18_mAd556_2 CB@18_mAd557_1 CB@18_mAd557_2 CB@18_mAd560_1 CB@18_mAd560_2 CB@18_mAd561_1 CB@18_mAd561_2 CB@18_mAd562_1 CB@18_mAd562_2 CB@18_mAd563_1 CB@18_mAd563_2 CB@18_mAd564_1 CB@18_mAd564_2 CB@18_mAd565_1 CB@18_mAd565_2 CB@18_mAd566_1 
+CB@18_mAd566_2 CB@18_mAd567_1 CB@18_mAd567_2 CB@18_mAd570_1 CB@18_mAd570_2 CB@18_mAd571_1 CB@18_mAd571_2 CB@18_mAd572_1 CB@18_mAd572_2 CB@18_mAd573_1 CB@18_mAd573_2 CB@18_mAd575_1 CB@18_mAd575_2 CB@18_mAd576_1 CB@18_mAd576_2 CB@18_mAd577_1 CB@18_mAd577_2 CB@18_mAd600_1 CB@18_mAd600_2 CB@18_mAd601_1 CB@18_mAd601_2 CB@18_mAd602_1 CB@18_mAd602_2 CB@18_mAd604_1 CB@18_mAd604_2 CB@18_mAd605_1 CB@18_mAd605_2 CB@18_mAd606_1 CB@18_mAd606_2 CB@18_mAd607_1 CB@18_mAd607_2 CB@18_mAd610_1 CB@18_mAd610_2 CB@18_mAd611_1 
+CB@18_mAd611_2 CB@18_mAd612_1 CB@18_mAd612_2 CB@18_mAd613_1 CB@18_mAd613_2 CB@18_mAd614_1 CB@18_mAd614_2 CB@18_mAd615_1 CB@18_mAd615_2 CB@18_mAd616_1 CB@18_mAd616_2 CB@18_mAd617_1 CB@18_mAd617_2 CB@18_mAd620_1 CB@18_mAd620_2 CB@18_mAd621_1 CB@18_mAd621_2 CB@18_mAd622_1 CB@18_mAd622_2 CB@18_mAd623_1 CB@18_mAd623_2 CB@18_mAd624_1 CB@18_mAd624_2 CB@18_mAd625_1 CB@18_mAd625_2 CB@18_mAd626_1 CB@18_mAd626_2 CB@18_mAd627_1 CB@18_mAd627_2 CB@18_mAd630_1 CB@18_mAd630_2 CB@18_mAd631_1 CB@18_mAd631_2 CB@18_mAd632_1 
+CB@18_mAd632_2 CB@18_mAd633_1 CB@18_mAd633_2 CB@18_mAd634_1 CB@18_mAd634_2 CB@18_mAd635_1 CB@18_mAd635_2 CB@18_mAd636_1 CB@18_mAd636_2 CB@18_mAd637_1 CB@18_mAd637_2 CB@18_mAd640_1 CB@18_mAd640_2 CB@18_mAd641_1 CB@18_mAd641_2 CB@18_mAd642_1 CB@18_mAd642_2 CB@18_mAd643_1 CB@18_mAd643_2 CB@18_mAd644_1 CB@18_mAd644_2 CB@18_mAd645_1 CB@18_mAd645_2 CB@18_mAd646_1 CB@18_mAd646_2 CB@18_mAd647_1 CB@18_mAd647_2 CB@18_mAd650_1 CB@18_mAd650_2 CB@18_mAd651_1 CB@18_mAd651_2 CB@18_mAd652_1 CB@18_mAd652_2 CB@18_mAd653_1 
+CB@18_mAd653_2 CB@18_mAd654_1 CB@18_mAd654_2 CB@18_mAd655_1 CB@18_mAd655_2 CB@18_mAd656_1 CB@18_mAd656_2 CB@18_mAd657_1 CB@18_mAd657_2 CB@18_mAd660_1 CB@18_mAd660_2 CB@18_mAd661_1 CB@18_mAd661_2 CB@18_mAd662_1 CB@18_mAd662_2 CB@18_mAd663_1 CB@18_mAd663_2 CB@18_mAd664_1 CB@18_mAd664_2 CB@18_mAd665_1 CB@18_mAd665_2 CB@18_mAd666_1 CB@18_mAd666_2 CB@18_mAd667_1 CB@18_mAd667_2 CB@18_mAd675_1 CB@18_mAd675_2 CB@18_mAd676_1 CB@18_mAd676_2 CB@18_mAd677_1 CB@18_mAd677_2 CB@18_mAd700_1 CB@18_mAd700_2 CB@18_mAd710_1 
+CB@18_mAd710_2 CB@18_mAd711_1 CB@18_mAd711_2 CB@18_mAd717_1 CB@18_mAd717_2 CB@18_mAd720_1 CB@18_mAd720_2 CB@18_mAd721_1 CB@18_mAd721_2 CB@18_mAd722_1 CB@18_mAd722_2 CB@18_mAd723_1 CB@18_mAd723_2 CB@18_mAd724_1 CB@18_mAd724_2 CB@18_mAd725_1 CB@18_mAd725_2 CB@18_mAd726_1 CB@18_mAd726_2 CB@18_mAd727_1 CB@18_mAd727_2 CB@18_mAd730_1 CB@18_mAd730_2 CB@18_mAd731_1 CB@18_mAd731_2 CB@18_mAd732_1 CB@18_mAd732_2 CB@18_mAd733_1 CB@18_mAd733_2 CB@18_mAd734_1 CB@18_mAd734_2 CB@18_mAd735_1 CB@18_mAd735_2 CB@18_mAd736_1 
+CB@18_mAd736_2 CB@18_mAd737_1 CB@18_mAd737_2 CB@18_mAd740_1 CB@18_mAd740_2 CB@18_mAd741_1 CB@18_mAd741_2 CB@18_mAd742_1 CB@18_mAd742_2 CB@18_mAd743_1 CB@18_mAd743_2 CB@18_mAd744_1 CB@18_mAd744_2 CB@18_mAd745_1 CB@18_mAd745_2 CB@18_mAd746_1 CB@18_mAd746_2 CB@18_mAd747_1 CB@18_mAd747_2 CB@18_mAd750_1 CB@18_mAd750_2 CB@18_mAd751_1 CB@18_mAd751_2 CB@18_mAd752_1 CB@18_mAd752_2 CB@18_mAd753_1 CB@18_mAd753_2 CB@18_mAd754_1 CB@18_mAd754_2 CB@18_mAd755_1 CB@18_mAd755_2 CB@18_mAd756_1 CB@18_mAd756_2 CB@18_mAd757_1 
+CB@18_mAd757_2 CB@18_mAd760_1 CB@18_mAd760_2 CB@18_mAd761_1 CB@18_mAd761_2 CB@18_mAd762_1 CB@18_mAd762_2 CB@18_mAd763_1 CB@18_mAd763_2 CB@18_mAd764_1 CB@18_mAd764_2 CB@18_mAd765_1 CB@18_mAd765_2 CB@18_mAd766_1 CB@18_mAd766_2 CB@18_mAd767_1 CB@18_mAd767_2 CB@18_mAd771_1 CB@18_mAd771_2 CB@18_mAd772_1 CB@18_mAd772_2 CB@18_mAd773_1 CB@18_mAd773_2 CB@18_mAd774_1 CB@18_mAd774_2 CB@18_mAd775_1 CB@18_mAd775_2 CB@18_mAd776_1 CB@18_mAd776_2 CB@18_mAd777_1 CB@18_mAd777_2 CB@18_X0 CB@18_X1 CB@18_X10 CB@18_X11 
+CB@18_X12 CB@18_X13 CB@18_X2 CB@18_X3 CB@18_X4 CB@18_X5 CB@18_X6 CB@18_X7 CB@18_X8 CB@18_X9 CB@18_Y1 CB@18_Y10 CB@18_Y11 CB@18_Y12 CB@18_Y2 CB@18_Y3 CB@18_Y4 CB@18_Y5 CB@18_Y6 CB@18_Y7 CB@18_Y8 CB@18_Y9 CB@18_Z1 CB@18_Z10 CB@18_Z11 CB@18_Z12 CB@18_Z2 CB@18_Z3 CB@18_Z4 CB@18_Z5 CB@18_Z6 CB@18_Z7 CB@18_Z8 CB@18_Z9 _5400TP094__CB
XCB@19 CB@19_K0 CB@19_K1 CB@19_K10 CB@19_K11 CB@19_K12 CB@19_K13 CB@19_K2 CB@19_K3 CB@19_K4 CB@19_K5 CB@19_K6 CB@19_K7 CB@19_K8 CB@19_K9 CB@19_mAd000_1 CB@19_mAd000_2 CB@19_mAd001_1 CB@19_mAd001_2 CB@19_mAd002_1 CB@19_mAd002_2 CB@19_mAd003_1 CB@19_mAd003_2 CB@19_mAd004_1 CB@19_mAd004_2 CB@19_mAd005_1 CB@19_mAd005_2 CB@19_mAd006_1 CB@19_mAd006_2 CB@19_mAd007_1 CB@19_mAd007_2 CB@19_mAd010_1 CB@19_mAd010_2 CB@19_mAd011_1 CB@19_mAd011_2 CB@19_mAd012_1 CB@19_mAd012_2 CB@19_mAd013_1 CB@19_mAd013_2 CB@19_mAd014_1 
+CB@19_mAd014_2 CB@19_mAd015_1 CB@19_mAd015_2 CB@19_mAd016_1 CB@19_mAd016_2 CB@19_mAd017_1 CB@19_mAd017_2 CB@19_mAd020_1 CB@19_mAd020_2 CB@19_mAd021_1 CB@19_mAd021_2 CB@19_mAd022_1 CB@19_mAd022_2 CB@19_mAd023_1 CB@19_mAd023_2 CB@19_mAd024_1 CB@19_mAd024_2 CB@19_mAd025_1 CB@19_mAd025_2 CB@19_mAd026_1 CB@19_mAd026_2 CB@19_mAd027_1 CB@19_mAd027_2 CB@19_mAd030_1 CB@19_mAd030_2 CB@19_mAd031_1 CB@19_mAd031_2 CB@19_mAd032_1 CB@19_mAd032_2 CB@19_mAd033_1 CB@19_mAd033_2 CB@19_mAd034_1 CB@19_mAd034_2 CB@19_mAd035_1 
+CB@19_mAd035_2 CB@19_mAd036_1 CB@19_mAd036_2 CB@19_mAd037_1 CB@19_mAd037_2 CB@19_mAd040_1 CB@19_mAd040_2 CB@19_mAd041_1 CB@19_mAd041_2 CB@19_mAd042_1 CB@19_mAd042_2 CB@19_mAd043_1 CB@19_mAd043_2 CB@19_mAd044_1 CB@19_mAd044_2 CB@19_mAd045_1 CB@19_mAd045_2 CB@19_mAd046_1 CB@19_mAd046_2 CB@19_mAd047_1 CB@19_mAd047_2 CB@19_mAd050_1 CB@19_mAd050_2 CB@19_mAd051_1 CB@19_mAd051_2 CB@19_mAd052_1 CB@19_mAd052_2 CB@19_mAd053_1 CB@19_mAd053_2 CB@19_mAd054_1 CB@19_mAd054_2 CB@19_mAd055_1 CB@19_mAd055_2 CB@19_mAd056_1 
+CB@19_mAd056_2 CB@19_mAd057_1 CB@19_mAd057_2 CB@19_mAd060_1 CB@19_mAd060_2 CB@19_mAd066_1 CB@19_mAd066_2 CB@19_mAd067_1 CB@19_mAd067_2 CB@19_mAd100_1 CB@19_mAd100_2 CB@19_mAd101_1 CB@19_mAd101_2 CB@19_mAd102_1 CB@19_mAd102_2 CB@19_mAd110_1 CB@19_mAd110_2 CB@19_mAd111_1 CB@19_mAd111_2 CB@19_mAd112_1 CB@19_mAd112_2 CB@19_mAd113_1 CB@19_mAd113_2 CB@19_mAd114_1 CB@19_mAd114_2 CB@19_mAd115_1 CB@19_mAd115_2 CB@19_mAd116_1 CB@19_mAd116_2 CB@19_mAd117_1 CB@19_mAd117_2 CB@19_mAd120_1 CB@19_mAd120_2 CB@19_mAd121_1 
+CB@19_mAd121_2 CB@19_mAd122_1 CB@19_mAd122_2 CB@19_mAd123_1 CB@19_mAd123_2 CB@19_mAd124_1 CB@19_mAd124_2 CB@19_mAd125_1 CB@19_mAd125_2 CB@19_mAd126_1 CB@19_mAd126_2 CB@19_mAd127_1 CB@19_mAd127_2 CB@19_mAd130_1 CB@19_mAd130_2 CB@19_mAd131_1 CB@19_mAd131_2 CB@19_mAd132_1 CB@19_mAd132_2 CB@19_mAd133_1 CB@19_mAd133_2 CB@19_mAd134_1 CB@19_mAd134_2 CB@19_mAd135_1 CB@19_mAd135_2 CB@19_mAd136_1 CB@19_mAd136_2 CB@19_mAd137_1 CB@19_mAd137_2 CB@19_mAd140_1 CB@19_mAd140_2 CB@19_mAd141_1 CB@19_mAd141_2 CB@19_mAd142_1 
+CB@19_mAd142_2 CB@19_mAd143_1 CB@19_mAd143_2 CB@19_mAd144_1 CB@19_mAd144_2 CB@19_mAd145_1 CB@19_mAd145_2 CB@19_mAd146_1 CB@19_mAd146_2 CB@19_mAd147_1 CB@19_mAd147_2 CB@19_mAd150_1 CB@19_mAd150_2 CB@19_mAd151_1 CB@19_mAd151_2 CB@19_mAd152_1 CB@19_mAd152_2 CB@19_mAd153_1 CB@19_mAd153_2 CB@19_mAd154_1 CB@19_mAd154_2 CB@19_mAd155_1 CB@19_mAd155_2 CB@19_mAd156_1 CB@19_mAd156_2 CB@19_mAd157_1 CB@19_mAd157_2 CB@19_mAd160_1 CB@19_mAd160_2 CB@19_mAd161_1 CB@19_mAd161_2 CB@19_mAd162_1 CB@19_mAd162_2 CB@19_mAd163_1 
+CB@19_mAd163_2 CB@19_mAd164_1 CB@19_mAd164_2 CB@19_mAd165_1 CB@19_mAd165_2 CB@19_mAd166_1 CB@19_mAd166_2 CB@19_mAd167_1 CB@19_mAd167_2 CB@19_mAd170_1 CB@19_mAd170_2 CB@19_mAd171_1 CB@19_mAd171_2 CB@19_mAd172_1 CB@19_mAd172_2 CB@19_mAd173_1 CB@19_mAd173_2 CB@19_mAd175_1 CB@19_mAd175_2 CB@19_mAd176_1 CB@19_mAd176_2 CB@19_mAd177_1 CB@19_mAd177_2 CB@19_mAd200_1 CB@19_mAd200_2 CB@19_mAd201_1 CB@19_mAd201_2 CB@19_mAd202_1 CB@19_mAd202_2 CB@19_mAd204_1 CB@19_mAd204_2 CB@19_mAd205_1 CB@19_mAd205_2 CB@19_mAd206_1 
+CB@19_mAd206_2 CB@19_mAd207_1 CB@19_mAd207_2 CB@19_mAd210_1 CB@19_mAd210_2 CB@19_mAd211_1 CB@19_mAd211_2 CB@19_mAd212_1 CB@19_mAd212_2 CB@19_mAd213_1 CB@19_mAd213_2 CB@19_mAd214_1 CB@19_mAd214_2 CB@19_mAd215_1 CB@19_mAd215_2 CB@19_mAd216_1 CB@19_mAd216_2 CB@19_mAd217_1 CB@19_mAd217_2 CB@19_mAd220_1 CB@19_mAd220_2 CB@19_mAd221_1 CB@19_mAd221_2 CB@19_mAd222_1 CB@19_mAd222_2 CB@19_mAd223_1 CB@19_mAd223_2 CB@19_mAd224_1 CB@19_mAd224_2 CB@19_mAd225_1 CB@19_mAd225_2 CB@19_mAd226_1 CB@19_mAd226_2 CB@19_mAd227_1 
+CB@19_mAd227_2 CB@19_mAd230_1 CB@19_mAd230_2 CB@19_mAd231_1 CB@19_mAd231_2 CB@19_mAd232_1 CB@19_mAd232_2 CB@19_mAd233_1 CB@19_mAd233_2 CB@19_mAd234_1 CB@19_mAd234_2 CB@19_mAd235_1 CB@19_mAd235_2 CB@19_mAd236_1 CB@19_mAd236_2 CB@19_mAd237_1 CB@19_mAd237_2 CB@19_mAd240_1 CB@19_mAd240_2 CB@19_mAd241_1 CB@19_mAd241_2 CB@19_mAd242_1 CB@19_mAd242_2 CB@19_mAd243_1 CB@19_mAd243_2 CB@19_mAd244_1 CB@19_mAd244_2 CB@19_mAd245_1 CB@19_mAd245_2 CB@19_mAd246_1 CB@19_mAd246_2 CB@19_mAd247_1 CB@19_mAd247_2 CB@19_mAd250_1 
+CB@19_mAd250_2 CB@19_mAd251_1 CB@19_mAd251_2 CB@19_mAd252_1 CB@19_mAd252_2 CB@19_mAd253_1 CB@19_mAd253_2 CB@19_mAd254_1 CB@19_mAd254_2 CB@19_mAd255_1 CB@19_mAd255_2 CB@19_mAd256_1 CB@19_mAd256_2 CB@19_mAd257_1 CB@19_mAd257_2 CB@19_mAd260_1 CB@19_mAd260_2 CB@19_mAd261_1 CB@19_mAd261_2 CB@19_mAd262_1 CB@19_mAd262_2 CB@19_mAd263_1 CB@19_mAd263_2 CB@19_mAd264_1 CB@19_mAd264_2 CB@19_mAd265_1 CB@19_mAd265_2 CB@19_mAd266_1 CB@19_mAd266_2 CB@19_mAd267_1 CB@19_mAd267_2 CB@19_mAd275_1 CB@19_mAd275_2 CB@19_mAd276_1 
+CB@19_mAd276_2 CB@19_mAd277_1 CB@19_mAd277_2 CB@19_mAd300_1 CB@19_mAd300_2 CB@19_mAd310_1 CB@19_mAd310_2 CB@19_mAd311_1 CB@19_mAd311_2 CB@19_mAd317_1 CB@19_mAd317_2 CB@19_mAd320_1 CB@19_mAd320_2 CB@19_mAd321_1 CB@19_mAd321_2 CB@19_mAd322_1 CB@19_mAd322_2 CB@19_mAd323_1 CB@19_mAd323_2 CB@19_mAd324_1 CB@19_mAd324_2 CB@19_mAd325_1 CB@19_mAd325_2 CB@19_mAd326_1 CB@19_mAd326_2 CB@19_mAd327_1 CB@19_mAd327_2 CB@19_mAd330_1 CB@19_mAd330_2 CB@19_mAd331_1 CB@19_mAd331_2 CB@19_mAd332_1 CB@19_mAd332_2 CB@19_mAd333_1 
+CB@19_mAd333_2 CB@19_mAd334_1 CB@19_mAd334_2 CB@19_mAd335_1 CB@19_mAd335_2 CB@19_mAd336_1 CB@19_mAd336_2 CB@19_mAd337_1 CB@19_mAd337_2 CB@19_mAd340_1 CB@19_mAd340_2 CB@19_mAd341_1 CB@19_mAd341_2 CB@19_mAd342_1 CB@19_mAd342_2 CB@19_mAd343_1 CB@19_mAd343_2 CB@19_mAd344_1 CB@19_mAd344_2 CB@19_mAd345_1 CB@19_mAd345_2 CB@19_mAd346_1 CB@19_mAd346_2 CB@19_mAd347_1 CB@19_mAd347_2 CB@19_mAd350_1 CB@19_mAd350_2 CB@19_mAd351_1 CB@19_mAd351_2 CB@19_mAd352_1 CB@19_mAd352_2 CB@19_mAd353_1 CB@19_mAd353_2 CB@19_mAd354_1 
+CB@19_mAd354_2 CB@19_mAd355_1 CB@19_mAd355_2 CB@19_mAd356_1 CB@19_mAd356_2 CB@19_mAd357_1 CB@19_mAd357_2 CB@19_mAd360_1 CB@19_mAd360_2 CB@19_mAd361_1 CB@19_mAd361_2 CB@19_mAd362_1 CB@19_mAd362_2 CB@19_mAd363_1 CB@19_mAd363_2 CB@19_mAd364_1 CB@19_mAd364_2 CB@19_mAd365_1 CB@19_mAd365_2 CB@19_mAd366_1 CB@19_mAd366_2 CB@19_mAd367_1 CB@19_mAd367_2 CB@19_mAd371_1 CB@19_mAd371_2 CB@19_mAd372_1 CB@19_mAd372_2 CB@19_mAd373_1 CB@19_mAd373_2 CB@19_mAd374_1 CB@19_mAd374_2 CB@19_mAd375_1 CB@19_mAd375_2 CB@19_mAd376_1 
+CB@19_mAd376_2 CB@19_mAd377_1 CB@19_mAd377_2 CB@19_mAd400_1 CB@19_mAd400_2 CB@19_mAd401_1 CB@19_mAd401_2 CB@19_mAd402_1 CB@19_mAd402_2 CB@19_mAd403_1 CB@19_mAd403_2 CB@19_mAd404_1 CB@19_mAd404_2 CB@19_mAd405_1 CB@19_mAd405_2 CB@19_mAd406_1 CB@19_mAd406_2 CB@19_mAd407_1 CB@19_mAd407_2 CB@19_mAd410_1 CB@19_mAd410_2 CB@19_mAd411_1 CB@19_mAd411_2 CB@19_mAd412_1 CB@19_mAd412_2 CB@19_mAd413_1 CB@19_mAd413_2 CB@19_mAd414_1 CB@19_mAd414_2 CB@19_mAd415_1 CB@19_mAd415_2 CB@19_mAd416_1 CB@19_mAd416_2 CB@19_mAd417_1 
+CB@19_mAd417_2 CB@19_mAd420_1 CB@19_mAd420_2 CB@19_mAd421_1 CB@19_mAd421_2 CB@19_mAd422_1 CB@19_mAd422_2 CB@19_mAd423_1 CB@19_mAd423_2 CB@19_mAd424_1 CB@19_mAd424_2 CB@19_mAd425_1 CB@19_mAd425_2 CB@19_mAd426_1 CB@19_mAd426_2 CB@19_mAd427_1 CB@19_mAd427_2 CB@19_mAd430_1 CB@19_mAd430_2 CB@19_mAd431_1 CB@19_mAd431_2 CB@19_mAd432_1 CB@19_mAd432_2 CB@19_mAd433_1 CB@19_mAd433_2 CB@19_mAd434_1 CB@19_mAd434_2 CB@19_mAd435_1 CB@19_mAd435_2 CB@19_mAd436_1 CB@19_mAd436_2 CB@19_mAd437_1 CB@19_mAd437_2 CB@19_mAd440_1 
+CB@19_mAd440_2 CB@19_mAd441_1 CB@19_mAd441_2 CB@19_mAd442_1 CB@19_mAd442_2 CB@19_mAd443_1 CB@19_mAd443_2 CB@19_mAd444_1 CB@19_mAd444_2 CB@19_mAd445_1 CB@19_mAd445_2 CB@19_mAd446_1 CB@19_mAd446_2 CB@19_mAd447_1 CB@19_mAd447_2 CB@19_mAd450_1 CB@19_mAd450_2 CB@19_mAd451_1 CB@19_mAd451_2 CB@19_mAd452_1 CB@19_mAd452_2 CB@19_mAd453_1 CB@19_mAd453_2 CB@19_mAd454_1 CB@19_mAd454_2 CB@19_mAd455_1 CB@19_mAd455_2 CB@19_mAd456_1 CB@19_mAd456_2 CB@19_mAd457_1 CB@19_mAd457_2 CB@19_mAd460_1 CB@19_mAd460_2 CB@19_mAd466_1 
+CB@19_mAd466_2 CB@19_mAd467_1 CB@19_mAd467_2 CB@19_mAd500_1 CB@19_mAd500_2 CB@19_mAd501_1 CB@19_mAd501_2 CB@19_mAd502_1 CB@19_mAd502_2 CB@19_mAd508_1 CB@19_mAd508_2 CB@19_mAd509_1 CB@19_mAd509_2 CB@19_mAd512_1 CB@19_mAd512_2 CB@19_mAd513_1 CB@19_mAd513_2 CB@19_mAd514_1 CB@19_mAd514_2 CB@19_mAd515_1 CB@19_mAd515_2 CB@19_mAd516_1 CB@19_mAd516_2 CB@19_mAd517_1 CB@19_mAd517_2 CB@19_mAd520_1 CB@19_mAd520_2 CB@19_mAd521_1 CB@19_mAd521_2 CB@19_mAd522_1 CB@19_mAd522_2 CB@19_mAd523_1 CB@19_mAd523_2 CB@19_mAd524_1 
+CB@19_mAd524_2 CB@19_mAd525_1 CB@19_mAd525_2 CB@19_mAd526_1 CB@19_mAd526_2 CB@19_mAd527_1 CB@19_mAd527_2 CB@19_mAd530_1 CB@19_mAd530_2 CB@19_mAd531_1 CB@19_mAd531_2 CB@19_mAd532_1 CB@19_mAd532_2 CB@19_mAd533_1 CB@19_mAd533_2 CB@19_mAd534_1 CB@19_mAd534_2 CB@19_mAd535_1 CB@19_mAd535_2 CB@19_mAd536_1 CB@19_mAd536_2 CB@19_mAd537_1 CB@19_mAd537_2 CB@19_mAd540_1 CB@19_mAd540_2 CB@19_mAd541_1 CB@19_mAd541_2 CB@19_mAd542_1 CB@19_mAd542_2 CB@19_mAd543_1 CB@19_mAd543_2 CB@19_mAd544_1 CB@19_mAd544_2 CB@19_mAd545_1 
+CB@19_mAd545_2 CB@19_mAd546_1 CB@19_mAd546_2 CB@19_mAd547_1 CB@19_mAd547_2 CB@19_mAd550_1 CB@19_mAd550_2 CB@19_mAd551_1 CB@19_mAd551_2 CB@19_mAd552_1 CB@19_mAd552_2 CB@19_mAd553_1 CB@19_mAd553_2 CB@19_mAd554_1 CB@19_mAd554_2 CB@19_mAd555_1 CB@19_mAd555_2 CB@19_mAd556_1 CB@19_mAd556_2 CB@19_mAd557_1 CB@19_mAd557_2 CB@19_mAd560_1 CB@19_mAd560_2 CB@19_mAd561_1 CB@19_mAd561_2 CB@19_mAd562_1 CB@19_mAd562_2 CB@19_mAd563_1 CB@19_mAd563_2 CB@19_mAd564_1 CB@19_mAd564_2 CB@19_mAd565_1 CB@19_mAd565_2 CB@19_mAd566_1 
+CB@19_mAd566_2 CB@19_mAd567_1 CB@19_mAd567_2 CB@19_mAd570_1 CB@19_mAd570_2 CB@19_mAd571_1 CB@19_mAd571_2 CB@19_mAd572_1 CB@19_mAd572_2 CB@19_mAd573_1 CB@19_mAd573_2 CB@19_mAd575_1 CB@19_mAd575_2 CB@19_mAd576_1 CB@19_mAd576_2 CB@19_mAd577_1 CB@19_mAd577_2 CB@19_mAd600_1 CB@19_mAd600_2 CB@19_mAd601_1 CB@19_mAd601_2 CB@19_mAd602_1 CB@19_mAd602_2 CB@19_mAd604_1 CB@19_mAd604_2 CB@19_mAd605_1 CB@19_mAd605_2 CB@19_mAd606_1 CB@19_mAd606_2 CB@19_mAd607_1 CB@19_mAd607_2 CB@19_mAd610_1 CB@19_mAd610_2 CB@19_mAd611_1 
+CB@19_mAd611_2 CB@19_mAd612_1 CB@19_mAd612_2 CB@19_mAd613_1 CB@19_mAd613_2 CB@19_mAd614_1 CB@19_mAd614_2 CB@19_mAd615_1 CB@19_mAd615_2 CB@19_mAd616_1 CB@19_mAd616_2 CB@19_mAd617_1 CB@19_mAd617_2 CB@19_mAd620_1 CB@19_mAd620_2 CB@19_mAd621_1 CB@19_mAd621_2 CB@19_mAd622_1 CB@19_mAd622_2 CB@19_mAd623_1 CB@19_mAd623_2 CB@19_mAd624_1 CB@19_mAd624_2 CB@19_mAd625_1 CB@19_mAd625_2 CB@19_mAd626_1 CB@19_mAd626_2 CB@19_mAd627_1 CB@19_mAd627_2 CB@19_mAd630_1 CB@19_mAd630_2 CB@19_mAd631_1 CB@19_mAd631_2 CB@19_mAd632_1 
+CB@19_mAd632_2 CB@19_mAd633_1 CB@19_mAd633_2 CB@19_mAd634_1 CB@19_mAd634_2 CB@19_mAd635_1 CB@19_mAd635_2 CB@19_mAd636_1 CB@19_mAd636_2 CB@19_mAd637_1 CB@19_mAd637_2 CB@19_mAd640_1 CB@19_mAd640_2 CB@19_mAd641_1 CB@19_mAd641_2 CB@19_mAd642_1 CB@19_mAd642_2 CB@19_mAd643_1 CB@19_mAd643_2 CB@19_mAd644_1 CB@19_mAd644_2 CB@19_mAd645_1 CB@19_mAd645_2 CB@19_mAd646_1 CB@19_mAd646_2 CB@19_mAd647_1 CB@19_mAd647_2 CB@19_mAd650_1 CB@19_mAd650_2 CB@19_mAd651_1 CB@19_mAd651_2 CB@19_mAd652_1 CB@19_mAd652_2 CB@19_mAd653_1 
+CB@19_mAd653_2 CB@19_mAd654_1 CB@19_mAd654_2 CB@19_mAd655_1 CB@19_mAd655_2 CB@19_mAd656_1 CB@19_mAd656_2 CB@19_mAd657_1 CB@19_mAd657_2 CB@19_mAd660_1 CB@19_mAd660_2 CB@19_mAd661_1 CB@19_mAd661_2 CB@19_mAd662_1 CB@19_mAd662_2 CB@19_mAd663_1 CB@19_mAd663_2 CB@19_mAd664_1 CB@19_mAd664_2 CB@19_mAd665_1 CB@19_mAd665_2 CB@19_mAd666_1 CB@19_mAd666_2 CB@19_mAd667_1 CB@19_mAd667_2 CB@19_mAd675_1 CB@19_mAd675_2 CB@19_mAd676_1 CB@19_mAd676_2 CB@19_mAd677_1 CB@19_mAd677_2 CB@19_mAd700_1 CB@19_mAd700_2 CB@19_mAd710_1 
+CB@19_mAd710_2 CB@19_mAd711_1 CB@19_mAd711_2 CB@19_mAd717_1 CB@19_mAd717_2 CB@19_mAd720_1 CB@19_mAd720_2 CB@19_mAd721_1 CB@19_mAd721_2 CB@19_mAd722_1 CB@19_mAd722_2 CB@19_mAd723_1 CB@19_mAd723_2 CB@19_mAd724_1 CB@19_mAd724_2 CB@19_mAd725_1 CB@19_mAd725_2 CB@19_mAd726_1 CB@19_mAd726_2 CB@19_mAd727_1 CB@19_mAd727_2 CB@19_mAd730_1 CB@19_mAd730_2 CB@19_mAd731_1 CB@19_mAd731_2 CB@19_mAd732_1 CB@19_mAd732_2 CB@19_mAd733_1 CB@19_mAd733_2 CB@19_mAd734_1 CB@19_mAd734_2 CB@19_mAd735_1 CB@19_mAd735_2 CB@19_mAd736_1 
+CB@19_mAd736_2 CB@19_mAd737_1 CB@19_mAd737_2 CB@19_mAd740_1 CB@19_mAd740_2 CB@19_mAd741_1 CB@19_mAd741_2 CB@19_mAd742_1 CB@19_mAd742_2 CB@19_mAd743_1 CB@19_mAd743_2 CB@19_mAd744_1 CB@19_mAd744_2 CB@19_mAd745_1 CB@19_mAd745_2 CB@19_mAd746_1 CB@19_mAd746_2 CB@19_mAd747_1 CB@19_mAd747_2 CB@19_mAd750_1 CB@19_mAd750_2 CB@19_mAd751_1 CB@19_mAd751_2 CB@19_mAd752_1 CB@19_mAd752_2 CB@19_mAd753_1 CB@19_mAd753_2 CB@19_mAd754_1 CB@19_mAd754_2 CB@19_mAd755_1 CB@19_mAd755_2 CB@19_mAd756_1 CB@19_mAd756_2 CB@19_mAd757_1 
+CB@19_mAd757_2 CB@19_mAd760_1 CB@19_mAd760_2 CB@19_mAd761_1 CB@19_mAd761_2 CB@19_mAd762_1 CB@19_mAd762_2 CB@19_mAd763_1 CB@19_mAd763_2 CB@19_mAd764_1 CB@19_mAd764_2 CB@19_mAd765_1 CB@19_mAd765_2 CB@19_mAd766_1 CB@19_mAd766_2 CB@19_mAd767_1 CB@19_mAd767_2 CB@19_mAd771_1 CB@19_mAd771_2 CB@19_mAd772_1 CB@19_mAd772_2 CB@19_mAd773_1 CB@19_mAd773_2 CB@19_mAd774_1 CB@19_mAd774_2 CB@19_mAd775_1 CB@19_mAd775_2 CB@19_mAd776_1 CB@19_mAd776_2 CB@19_mAd777_1 CB@19_mAd777_2 CB@19_X0 CB@19_X1 CB@19_X10 CB@19_X11 
+CB@19_X12 CB@19_X13 CB@19_X2 CB@19_X3 CB@19_X4 CB@19_X5 CB@19_X6 CB@19_X7 CB@19_X8 CB@19_X9 CB@19_Y1 CB@19_Y10 CB@19_Y11 CB@19_Y12 CB@19_Y2 CB@19_Y3 CB@19_Y4 CB@19_Y5 CB@19_Y6 CB@19_Y7 CB@19_Y8 CB@19_Y9 CB@19_Z1 CB@19_Z10 CB@19_Z11 CB@19_Z12 CB@19_Z2 CB@19_Z3 CB@19_Z4 CB@19_Z5 CB@19_Z6 CB@19_Z7 CB@19_Z8 CB@19_Z9 _5400TP094__CB
XCB@20 CB@20_K0 CB@20_K1 CB@20_K10 CB@20_K11 CB@20_K12 CB@20_K13 CB@20_K2 CB@20_K3 CB@20_K4 CB@20_K5 CB@20_K6 CB@20_K7 CB@20_K8 CB@20_K9 CB@20_mAd000_1 CB@20_mAd000_2 CB@20_mAd001_1 CB@20_mAd001_2 CB@20_mAd002_1 CB@20_mAd002_2 CB@20_mAd003_1 CB@20_mAd003_2 CB@20_mAd004_1 CB@20_mAd004_2 CB@20_mAd005_1 CB@20_mAd005_2 CB@20_mAd006_1 CB@20_mAd006_2 CB@20_mAd007_1 CB@20_mAd007_2 CB@20_mAd010_1 CB@20_mAd010_2 CB@20_mAd011_1 CB@20_mAd011_2 CB@20_mAd012_1 CB@20_mAd012_2 CB@20_mAd013_1 CB@20_mAd013_2 CB@20_mAd014_1 
+CB@20_mAd014_2 CB@20_mAd015_1 CB@20_mAd015_2 CB@20_mAd016_1 CB@20_mAd016_2 CB@20_mAd017_1 CB@20_mAd017_2 CB@20_mAd020_1 CB@20_mAd020_2 CB@20_mAd021_1 CB@20_mAd021_2 CB@20_mAd022_1 CB@20_mAd022_2 CB@20_mAd023_1 CB@20_mAd023_2 CB@20_mAd024_1 CB@20_mAd024_2 CB@20_mAd025_1 CB@20_mAd025_2 CB@20_mAd026_1 CB@20_mAd026_2 CB@20_mAd027_1 CB@20_mAd027_2 CB@20_mAd030_1 CB@20_mAd030_2 CB@20_mAd031_1 CB@20_mAd031_2 CB@20_mAd032_1 CB@20_mAd032_2 CB@20_mAd033_1 CB@20_mAd033_2 CB@20_mAd034_1 CB@20_mAd034_2 CB@20_mAd035_1 
+CB@20_mAd035_2 CB@20_mAd036_1 CB@20_mAd036_2 CB@20_mAd037_1 CB@20_mAd037_2 CB@20_mAd040_1 CB@20_mAd040_2 CB@20_mAd041_1 CB@20_mAd041_2 CB@20_mAd042_1 CB@20_mAd042_2 CB@20_mAd043_1 CB@20_mAd043_2 CB@20_mAd044_1 CB@20_mAd044_2 CB@20_mAd045_1 CB@20_mAd045_2 CB@20_mAd046_1 CB@20_mAd046_2 CB@20_mAd047_1 CB@20_mAd047_2 CB@20_mAd050_1 CB@20_mAd050_2 CB@20_mAd051_1 CB@20_mAd051_2 CB@20_mAd052_1 CB@20_mAd052_2 CB@20_mAd053_1 CB@20_mAd053_2 CB@20_mAd054_1 CB@20_mAd054_2 CB@20_mAd055_1 CB@20_mAd055_2 CB@20_mAd056_1 
+CB@20_mAd056_2 CB@20_mAd057_1 CB@20_mAd057_2 CB@20_mAd060_1 CB@20_mAd060_2 CB@20_mAd066_1 CB@20_mAd066_2 CB@20_mAd067_1 CB@20_mAd067_2 CB@20_mAd100_1 CB@20_mAd100_2 CB@20_mAd101_1 CB@20_mAd101_2 CB@20_mAd102_1 CB@20_mAd102_2 CB@20_mAd110_1 CB@20_mAd110_2 CB@20_mAd111_1 CB@20_mAd111_2 CB@20_mAd112_1 CB@20_mAd112_2 CB@20_mAd113_1 CB@20_mAd113_2 CB@20_mAd114_1 CB@20_mAd114_2 CB@20_mAd115_1 CB@20_mAd115_2 CB@20_mAd116_1 CB@20_mAd116_2 CB@20_mAd117_1 CB@20_mAd117_2 CB@20_mAd120_1 CB@20_mAd120_2 CB@20_mAd121_1 
+CB@20_mAd121_2 CB@20_mAd122_1 CB@20_mAd122_2 CB@20_mAd123_1 CB@20_mAd123_2 CB@20_mAd124_1 CB@20_mAd124_2 CB@20_mAd125_1 CB@20_mAd125_2 CB@20_mAd126_1 CB@20_mAd126_2 CB@20_mAd127_1 CB@20_mAd127_2 CB@20_mAd130_1 CB@20_mAd130_2 CB@20_mAd131_1 CB@20_mAd131_2 CB@20_mAd132_1 CB@20_mAd132_2 CB@20_mAd133_1 CB@20_mAd133_2 CB@20_mAd134_1 CB@20_mAd134_2 CB@20_mAd135_1 CB@20_mAd135_2 CB@20_mAd136_1 CB@20_mAd136_2 CB@20_mAd137_1 CB@20_mAd137_2 CB@20_mAd140_1 CB@20_mAd140_2 CB@20_mAd141_1 CB@20_mAd141_2 CB@20_mAd142_1 
+CB@20_mAd142_2 CB@20_mAd143_1 CB@20_mAd143_2 CB@20_mAd144_1 CB@20_mAd144_2 CB@20_mAd145_1 CB@20_mAd145_2 CB@20_mAd146_1 CB@20_mAd146_2 CB@20_mAd147_1 CB@20_mAd147_2 CB@20_mAd150_1 CB@20_mAd150_2 CB@20_mAd151_1 CB@20_mAd151_2 CB@20_mAd152_1 CB@20_mAd152_2 CB@20_mAd153_1 CB@20_mAd153_2 CB@20_mAd154_1 CB@20_mAd154_2 CB@20_mAd155_1 CB@20_mAd155_2 CB@20_mAd156_1 CB@20_mAd156_2 CB@20_mAd157_1 CB@20_mAd157_2 CB@20_mAd160_1 CB@20_mAd160_2 CB@20_mAd161_1 CB@20_mAd161_2 CB@20_mAd162_1 CB@20_mAd162_2 CB@20_mAd163_1 
+CB@20_mAd163_2 CB@20_mAd164_1 CB@20_mAd164_2 CB@20_mAd165_1 CB@20_mAd165_2 CB@20_mAd166_1 CB@20_mAd166_2 CB@20_mAd167_1 CB@20_mAd167_2 CB@20_mAd170_1 CB@20_mAd170_2 CB@20_mAd171_1 CB@20_mAd171_2 CB@20_mAd172_1 CB@20_mAd172_2 CB@20_mAd173_1 CB@20_mAd173_2 CB@20_mAd175_1 CB@20_mAd175_2 CB@20_mAd176_1 CB@20_mAd176_2 CB@20_mAd177_1 CB@20_mAd177_2 CB@20_mAd200_1 CB@20_mAd200_2 CB@20_mAd201_1 CB@20_mAd201_2 CB@20_mAd202_1 CB@20_mAd202_2 CB@20_mAd204_1 CB@20_mAd204_2 CB@20_mAd205_1 CB@20_mAd205_2 CB@20_mAd206_1 
+CB@20_mAd206_2 CB@20_mAd207_1 CB@20_mAd207_2 CB@20_mAd210_1 CB@20_mAd210_2 CB@20_mAd211_1 CB@20_mAd211_2 CB@20_mAd212_1 CB@20_mAd212_2 CB@20_mAd213_1 CB@20_mAd213_2 CB@20_mAd214_1 CB@20_mAd214_2 CB@20_mAd215_1 CB@20_mAd215_2 CB@20_mAd216_1 CB@20_mAd216_2 CB@20_mAd217_1 CB@20_mAd217_2 CB@20_mAd220_1 CB@20_mAd220_2 CB@20_mAd221_1 CB@20_mAd221_2 CB@20_mAd222_1 CB@20_mAd222_2 CB@20_mAd223_1 CB@20_mAd223_2 CB@20_mAd224_1 CB@20_mAd224_2 CB@20_mAd225_1 CB@20_mAd225_2 CB@20_mAd226_1 CB@20_mAd226_2 CB@20_mAd227_1 
+CB@20_mAd227_2 CB@20_mAd230_1 CB@20_mAd230_2 CB@20_mAd231_1 CB@20_mAd231_2 CB@20_mAd232_1 CB@20_mAd232_2 CB@20_mAd233_1 CB@20_mAd233_2 CB@20_mAd234_1 CB@20_mAd234_2 CB@20_mAd235_1 CB@20_mAd235_2 CB@20_mAd236_1 CB@20_mAd236_2 CB@20_mAd237_1 CB@20_mAd237_2 CB@20_mAd240_1 CB@20_mAd240_2 CB@20_mAd241_1 CB@20_mAd241_2 CB@20_mAd242_1 CB@20_mAd242_2 CB@20_mAd243_1 CB@20_mAd243_2 CB@20_mAd244_1 CB@20_mAd244_2 CB@20_mAd245_1 CB@20_mAd245_2 CB@20_mAd246_1 CB@20_mAd246_2 CB@20_mAd247_1 CB@20_mAd247_2 CB@20_mAd250_1 
+CB@20_mAd250_2 CB@20_mAd251_1 CB@20_mAd251_2 CB@20_mAd252_1 CB@20_mAd252_2 CB@20_mAd253_1 CB@20_mAd253_2 CB@20_mAd254_1 CB@20_mAd254_2 CB@20_mAd255_1 CB@20_mAd255_2 CB@20_mAd256_1 CB@20_mAd256_2 CB@20_mAd257_1 CB@20_mAd257_2 CB@20_mAd260_1 CB@20_mAd260_2 CB@20_mAd261_1 CB@20_mAd261_2 CB@20_mAd262_1 CB@20_mAd262_2 CB@20_mAd263_1 CB@20_mAd263_2 CB@20_mAd264_1 CB@20_mAd264_2 CB@20_mAd265_1 CB@20_mAd265_2 CB@20_mAd266_1 CB@20_mAd266_2 CB@20_mAd267_1 CB@20_mAd267_2 CB@20_mAd275_1 CB@20_mAd275_2 CB@20_mAd276_1 
+CB@20_mAd276_2 CB@20_mAd277_1 CB@20_mAd277_2 CB@20_mAd300_1 CB@20_mAd300_2 CB@20_mAd310_1 CB@20_mAd310_2 CB@20_mAd311_1 CB@20_mAd311_2 CB@20_mAd317_1 CB@20_mAd317_2 CB@20_mAd320_1 CB@20_mAd320_2 CB@20_mAd321_1 CB@20_mAd321_2 CB@20_mAd322_1 CB@20_mAd322_2 CB@20_mAd323_1 CB@20_mAd323_2 CB@20_mAd324_1 CB@20_mAd324_2 CB@20_mAd325_1 CB@20_mAd325_2 CB@20_mAd326_1 CB@20_mAd326_2 CB@20_mAd327_1 CB@20_mAd327_2 CB@20_mAd330_1 CB@20_mAd330_2 CB@20_mAd331_1 CB@20_mAd331_2 CB@20_mAd332_1 CB@20_mAd332_2 CB@20_mAd333_1 
+CB@20_mAd333_2 CB@20_mAd334_1 CB@20_mAd334_2 CB@20_mAd335_1 CB@20_mAd335_2 CB@20_mAd336_1 CB@20_mAd336_2 CB@20_mAd337_1 CB@20_mAd337_2 CB@20_mAd340_1 CB@20_mAd340_2 CB@20_mAd341_1 CB@20_mAd341_2 CB@20_mAd342_1 CB@20_mAd342_2 CB@20_mAd343_1 CB@20_mAd343_2 CB@20_mAd344_1 CB@20_mAd344_2 CB@20_mAd345_1 CB@20_mAd345_2 CB@20_mAd346_1 CB@20_mAd346_2 CB@20_mAd347_1 CB@20_mAd347_2 CB@20_mAd350_1 CB@20_mAd350_2 CB@20_mAd351_1 CB@20_mAd351_2 CB@20_mAd352_1 CB@20_mAd352_2 CB@20_mAd353_1 CB@20_mAd353_2 CB@20_mAd354_1 
+CB@20_mAd354_2 CB@20_mAd355_1 CB@20_mAd355_2 CB@20_mAd356_1 CB@20_mAd356_2 CB@20_mAd357_1 CB@20_mAd357_2 CB@20_mAd360_1 CB@20_mAd360_2 CB@20_mAd361_1 CB@20_mAd361_2 CB@20_mAd362_1 CB@20_mAd362_2 CB@20_mAd363_1 CB@20_mAd363_2 CB@20_mAd364_1 CB@20_mAd364_2 CB@20_mAd365_1 CB@20_mAd365_2 CB@20_mAd366_1 CB@20_mAd366_2 CB@20_mAd367_1 CB@20_mAd367_2 CB@20_mAd371_1 CB@20_mAd371_2 CB@20_mAd372_1 CB@20_mAd372_2 CB@20_mAd373_1 CB@20_mAd373_2 CB@20_mAd374_1 CB@20_mAd374_2 CB@20_mAd375_1 CB@20_mAd375_2 CB@20_mAd376_1 
+CB@20_mAd376_2 CB@20_mAd377_1 CB@20_mAd377_2 CB@20_mAd400_1 CB@20_mAd400_2 CB@20_mAd401_1 CB@20_mAd401_2 CB@20_mAd402_1 CB@20_mAd402_2 CB@20_mAd403_1 CB@20_mAd403_2 CB@20_mAd404_1 CB@20_mAd404_2 CB@20_mAd405_1 CB@20_mAd405_2 CB@20_mAd406_1 CB@20_mAd406_2 CB@20_mAd407_1 CB@20_mAd407_2 CB@20_mAd410_1 CB@20_mAd410_2 CB@20_mAd411_1 CB@20_mAd411_2 CB@20_mAd412_1 CB@20_mAd412_2 CB@20_mAd413_1 CB@20_mAd413_2 CB@20_mAd414_1 CB@20_mAd414_2 CB@20_mAd415_1 CB@20_mAd415_2 CB@20_mAd416_1 CB@20_mAd416_2 CB@20_mAd417_1 
+CB@20_mAd417_2 CB@20_mAd420_1 CB@20_mAd420_2 CB@20_mAd421_1 CB@20_mAd421_2 CB@20_mAd422_1 CB@20_mAd422_2 CB@20_mAd423_1 CB@20_mAd423_2 CB@20_mAd424_1 CB@20_mAd424_2 CB@20_mAd425_1 CB@20_mAd425_2 CB@20_mAd426_1 CB@20_mAd426_2 CB@20_mAd427_1 CB@20_mAd427_2 CB@20_mAd430_1 CB@20_mAd430_2 CB@20_mAd431_1 CB@20_mAd431_2 CB@20_mAd432_1 CB@20_mAd432_2 CB@20_mAd433_1 CB@20_mAd433_2 CB@20_mAd434_1 CB@20_mAd434_2 CB@20_mAd435_1 CB@20_mAd435_2 CB@20_mAd436_1 CB@20_mAd436_2 CB@20_mAd437_1 CB@20_mAd437_2 CB@20_mAd440_1 
+CB@20_mAd440_2 CB@20_mAd441_1 CB@20_mAd441_2 CB@20_mAd442_1 CB@20_mAd442_2 CB@20_mAd443_1 CB@20_mAd443_2 CB@20_mAd444_1 CB@20_mAd444_2 CB@20_mAd445_1 CB@20_mAd445_2 CB@20_mAd446_1 CB@20_mAd446_2 CB@20_mAd447_1 CB@20_mAd447_2 CB@20_mAd450_1 CB@20_mAd450_2 CB@20_mAd451_1 CB@20_mAd451_2 CB@20_mAd452_1 CB@20_mAd452_2 CB@20_mAd453_1 CB@20_mAd453_2 CB@20_mAd454_1 CB@20_mAd454_2 CB@20_mAd455_1 CB@20_mAd455_2 CB@20_mAd456_1 CB@20_mAd456_2 CB@20_mAd457_1 CB@20_mAd457_2 CB@20_mAd460_1 CB@20_mAd460_2 CB@20_mAd466_1 
+CB@20_mAd466_2 CB@20_mAd467_1 CB@20_mAd467_2 CB@20_mAd500_1 CB@20_mAd500_2 CB@20_mAd501_1 CB@20_mAd501_2 CB@20_mAd502_1 CB@20_mAd502_2 CB@20_mAd508_1 CB@20_mAd508_2 CB@20_mAd509_1 CB@20_mAd509_2 CB@20_mAd512_1 CB@20_mAd512_2 CB@20_mAd513_1 CB@20_mAd513_2 CB@20_mAd514_1 CB@20_mAd514_2 CB@20_mAd515_1 CB@20_mAd515_2 CB@20_mAd516_1 CB@20_mAd516_2 CB@20_mAd517_1 CB@20_mAd517_2 CB@20_mAd520_1 CB@20_mAd520_2 CB@20_mAd521_1 CB@20_mAd521_2 CB@20_mAd522_1 CB@20_mAd522_2 CB@20_mAd523_1 CB@20_mAd523_2 CB@20_mAd524_1 
+CB@20_mAd524_2 CB@20_mAd525_1 CB@20_mAd525_2 CB@20_mAd526_1 CB@20_mAd526_2 CB@20_mAd527_1 CB@20_mAd527_2 CB@20_mAd530_1 CB@20_mAd530_2 CB@20_mAd531_1 CB@20_mAd531_2 CB@20_mAd532_1 CB@20_mAd532_2 CB@20_mAd533_1 CB@20_mAd533_2 CB@20_mAd534_1 CB@20_mAd534_2 CB@20_mAd535_1 CB@20_mAd535_2 CB@20_mAd536_1 CB@20_mAd536_2 CB@20_mAd537_1 CB@20_mAd537_2 CB@20_mAd540_1 CB@20_mAd540_2 CB@20_mAd541_1 CB@20_mAd541_2 CB@20_mAd542_1 CB@20_mAd542_2 CB@20_mAd543_1 CB@20_mAd543_2 CB@20_mAd544_1 CB@20_mAd544_2 CB@20_mAd545_1 
+CB@20_mAd545_2 CB@20_mAd546_1 CB@20_mAd546_2 CB@20_mAd547_1 CB@20_mAd547_2 CB@20_mAd550_1 CB@20_mAd550_2 CB@20_mAd551_1 CB@20_mAd551_2 CB@20_mAd552_1 CB@20_mAd552_2 CB@20_mAd553_1 CB@20_mAd553_2 CB@20_mAd554_1 CB@20_mAd554_2 CB@20_mAd555_1 CB@20_mAd555_2 CB@20_mAd556_1 CB@20_mAd556_2 CB@20_mAd557_1 CB@20_mAd557_2 CB@20_mAd560_1 CB@20_mAd560_2 CB@20_mAd561_1 CB@20_mAd561_2 CB@20_mAd562_1 CB@20_mAd562_2 CB@20_mAd563_1 CB@20_mAd563_2 CB@20_mAd564_1 CB@20_mAd564_2 CB@20_mAd565_1 CB@20_mAd565_2 CB@20_mAd566_1 
+CB@20_mAd566_2 CB@20_mAd567_1 CB@20_mAd567_2 CB@20_mAd570_1 CB@20_mAd570_2 CB@20_mAd571_1 CB@20_mAd571_2 CB@20_mAd572_1 CB@20_mAd572_2 CB@20_mAd573_1 CB@20_mAd573_2 CB@20_mAd575_1 CB@20_mAd575_2 CB@20_mAd576_1 CB@20_mAd576_2 CB@20_mAd577_1 CB@20_mAd577_2 CB@20_mAd600_1 CB@20_mAd600_2 CB@20_mAd601_1 CB@20_mAd601_2 CB@20_mAd602_1 CB@20_mAd602_2 CB@20_mAd604_1 CB@20_mAd604_2 CB@20_mAd605_1 CB@20_mAd605_2 CB@20_mAd606_1 CB@20_mAd606_2 CB@20_mAd607_1 CB@20_mAd607_2 CB@20_mAd610_1 CB@20_mAd610_2 CB@20_mAd611_1 
+CB@20_mAd611_2 CB@20_mAd612_1 CB@20_mAd612_2 CB@20_mAd613_1 CB@20_mAd613_2 CB@20_mAd614_1 CB@20_mAd614_2 CB@20_mAd615_1 CB@20_mAd615_2 CB@20_mAd616_1 CB@20_mAd616_2 CB@20_mAd617_1 CB@20_mAd617_2 CB@20_mAd620_1 CB@20_mAd620_2 CB@20_mAd621_1 CB@20_mAd621_2 CB@20_mAd622_1 CB@20_mAd622_2 CB@20_mAd623_1 CB@20_mAd623_2 CB@20_mAd624_1 CB@20_mAd624_2 CB@20_mAd625_1 CB@20_mAd625_2 CB@20_mAd626_1 CB@20_mAd626_2 CB@20_mAd627_1 CB@20_mAd627_2 CB@20_mAd630_1 CB@20_mAd630_2 CB@20_mAd631_1 CB@20_mAd631_2 CB@20_mAd632_1 
+CB@20_mAd632_2 CB@20_mAd633_1 CB@20_mAd633_2 CB@20_mAd634_1 CB@20_mAd634_2 CB@20_mAd635_1 CB@20_mAd635_2 CB@20_mAd636_1 CB@20_mAd636_2 CB@20_mAd637_1 CB@20_mAd637_2 CB@20_mAd640_1 CB@20_mAd640_2 CB@20_mAd641_1 CB@20_mAd641_2 CB@20_mAd642_1 CB@20_mAd642_2 CB@20_mAd643_1 CB@20_mAd643_2 CB@20_mAd644_1 CB@20_mAd644_2 CB@20_mAd645_1 CB@20_mAd645_2 CB@20_mAd646_1 CB@20_mAd646_2 CB@20_mAd647_1 CB@20_mAd647_2 CB@20_mAd650_1 CB@20_mAd650_2 CB@20_mAd651_1 CB@20_mAd651_2 CB@20_mAd652_1 CB@20_mAd652_2 CB@20_mAd653_1 
+CB@20_mAd653_2 CB@20_mAd654_1 CB@20_mAd654_2 CB@20_mAd655_1 CB@20_mAd655_2 CB@20_mAd656_1 CB@20_mAd656_2 CB@20_mAd657_1 CB@20_mAd657_2 CB@20_mAd660_1 CB@20_mAd660_2 CB@20_mAd661_1 CB@20_mAd661_2 CB@20_mAd662_1 CB@20_mAd662_2 CB@20_mAd663_1 CB@20_mAd663_2 CB@20_mAd664_1 CB@20_mAd664_2 CB@20_mAd665_1 CB@20_mAd665_2 CB@20_mAd666_1 CB@20_mAd666_2 CB@20_mAd667_1 CB@20_mAd667_2 CB@20_mAd675_1 CB@20_mAd675_2 CB@20_mAd676_1 CB@20_mAd676_2 CB@20_mAd677_1 CB@20_mAd677_2 CB@20_mAd700_1 CB@20_mAd700_2 CB@20_mAd710_1 
+CB@20_mAd710_2 CB@20_mAd711_1 CB@20_mAd711_2 CB@20_mAd717_1 CB@20_mAd717_2 CB@20_mAd720_1 CB@20_mAd720_2 CB@20_mAd721_1 CB@20_mAd721_2 CB@20_mAd722_1 CB@20_mAd722_2 CB@20_mAd723_1 CB@20_mAd723_2 CB@20_mAd724_1 CB@20_mAd724_2 CB@20_mAd725_1 CB@20_mAd725_2 CB@20_mAd726_1 CB@20_mAd726_2 CB@20_mAd727_1 CB@20_mAd727_2 CB@20_mAd730_1 CB@20_mAd730_2 CB@20_mAd731_1 CB@20_mAd731_2 CB@20_mAd732_1 CB@20_mAd732_2 CB@20_mAd733_1 CB@20_mAd733_2 CB@20_mAd734_1 CB@20_mAd734_2 CB@20_mAd735_1 CB@20_mAd735_2 CB@20_mAd736_1 
+CB@20_mAd736_2 CB@20_mAd737_1 CB@20_mAd737_2 CB@20_mAd740_1 CB@20_mAd740_2 CB@20_mAd741_1 CB@20_mAd741_2 CB@20_mAd742_1 CB@20_mAd742_2 CB@20_mAd743_1 CB@20_mAd743_2 CB@20_mAd744_1 CB@20_mAd744_2 CB@20_mAd745_1 CB@20_mAd745_2 CB@20_mAd746_1 CB@20_mAd746_2 CB@20_mAd747_1 CB@20_mAd747_2 CB@20_mAd750_1 CB@20_mAd750_2 CB@20_mAd751_1 CB@20_mAd751_2 CB@20_mAd752_1 CB@20_mAd752_2 CB@20_mAd753_1 CB@20_mAd753_2 CB@20_mAd754_1 CB@20_mAd754_2 CB@20_mAd755_1 CB@20_mAd755_2 CB@20_mAd756_1 CB@20_mAd756_2 CB@20_mAd757_1 
+CB@20_mAd757_2 CB@20_mAd760_1 CB@20_mAd760_2 CB@20_mAd761_1 CB@20_mAd761_2 CB@20_mAd762_1 CB@20_mAd762_2 CB@20_mAd763_1 CB@20_mAd763_2 CB@20_mAd764_1 CB@20_mAd764_2 CB@20_mAd765_1 CB@20_mAd765_2 CB@20_mAd766_1 CB@20_mAd766_2 CB@20_mAd767_1 CB@20_mAd767_2 CB@20_mAd771_1 CB@20_mAd771_2 CB@20_mAd772_1 CB@20_mAd772_2 CB@20_mAd773_1 CB@20_mAd773_2 CB@20_mAd774_1 CB@20_mAd774_2 CB@20_mAd775_1 CB@20_mAd775_2 CB@20_mAd776_1 CB@20_mAd776_2 CB@20_mAd777_1 CB@20_mAd777_2 CB@20_X0 CB@20_X1 CB@20_X10 CB@20_X11 
+CB@20_X12 CB@20_X13 CB@20_X2 CB@20_X3 CB@20_X4 CB@20_X5 CB@20_X6 CB@20_X7 CB@20_X8 CB@20_X9 CB@20_Y1 CB@20_Y10 CB@20_Y11 CB@20_Y12 CB@20_Y2 CB@20_Y3 CB@20_Y4 CB@20_Y5 CB@20_Y6 CB@20_Y7 CB@20_Y8 CB@20_Y9 CB@20_Z1 CB@20_Z10 CB@20_Z11 CB@20_Z12 CB@20_Z2 CB@20_Z3 CB@20_Z4 CB@20_Z5 CB@20_Z6 CB@20_Z7 CB@20_Z8 CB@20_Z9 _5400TP094__CB
XCB@21 CB@21_K0 CB@21_K1 CB@21_K10 CB@21_K11 CB@21_K12 CB@21_K13 CB@21_K2 CB@21_K3 CB@21_K4 CB@21_K5 CB@21_K6 CB@21_K7 CB@21_K8 CB@21_K9 CB@21_mAd000_1 CB@21_mAd000_2 CB@21_mAd001_1 CB@21_mAd001_2 CB@21_mAd002_1 CB@21_mAd002_2 CB@21_mAd003_1 CB@21_mAd003_2 CB@21_mAd004_1 CB@21_mAd004_2 CB@21_mAd005_1 CB@21_mAd005_2 CB@21_mAd006_1 CB@21_mAd006_2 CB@21_mAd007_1 CB@21_mAd007_2 CB@21_mAd010_1 CB@21_mAd010_2 CB@21_mAd011_1 CB@21_mAd011_2 CB@21_mAd012_1 CB@21_mAd012_2 CB@21_mAd013_1 CB@21_mAd013_2 CB@21_mAd014_1 
+CB@21_mAd014_2 CB@21_mAd015_1 CB@21_mAd015_2 CB@21_mAd016_1 CB@21_mAd016_2 CB@21_mAd017_1 CB@21_mAd017_2 CB@21_mAd020_1 CB@21_mAd020_2 CB@21_mAd021_1 CB@21_mAd021_2 CB@21_mAd022_1 CB@21_mAd022_2 CB@21_mAd023_1 CB@21_mAd023_2 CB@21_mAd024_1 CB@21_mAd024_2 CB@21_mAd025_1 CB@21_mAd025_2 CB@21_mAd026_1 CB@21_mAd026_2 CB@21_mAd027_1 CB@21_mAd027_2 CB@21_mAd030_1 CB@21_mAd030_2 CB@21_mAd031_1 CB@21_mAd031_2 CB@21_mAd032_1 CB@21_mAd032_2 CB@21_mAd033_1 CB@21_mAd033_2 CB@21_mAd034_1 CB@21_mAd034_2 CB@21_mAd035_1 
+CB@21_mAd035_2 CB@21_mAd036_1 CB@21_mAd036_2 CB@21_mAd037_1 CB@21_mAd037_2 CB@21_mAd040_1 CB@21_mAd040_2 CB@21_mAd041_1 CB@21_mAd041_2 CB@21_mAd042_1 CB@21_mAd042_2 CB@21_mAd043_1 CB@21_mAd043_2 CB@21_mAd044_1 CB@21_mAd044_2 CB@21_mAd045_1 CB@21_mAd045_2 CB@21_mAd046_1 CB@21_mAd046_2 CB@21_mAd047_1 CB@21_mAd047_2 CB@21_mAd050_1 CB@21_mAd050_2 CB@21_mAd051_1 CB@21_mAd051_2 CB@21_mAd052_1 CB@21_mAd052_2 CB@21_mAd053_1 CB@21_mAd053_2 CB@21_mAd054_1 CB@21_mAd054_2 CB@21_mAd055_1 CB@21_mAd055_2 CB@21_mAd056_1 
+CB@21_mAd056_2 CB@21_mAd057_1 CB@21_mAd057_2 CB@21_mAd060_1 CB@21_mAd060_2 CB@21_mAd066_1 CB@21_mAd066_2 CB@21_mAd067_1 CB@21_mAd067_2 CB@21_mAd100_1 CB@21_mAd100_2 CB@21_mAd101_1 CB@21_mAd101_2 CB@21_mAd102_1 CB@21_mAd102_2 CB@21_mAd110_1 CB@21_mAd110_2 CB@21_mAd111_1 CB@21_mAd111_2 CB@21_mAd112_1 CB@21_mAd112_2 CB@21_mAd113_1 CB@21_mAd113_2 CB@21_mAd114_1 CB@21_mAd114_2 CB@21_mAd115_1 CB@21_mAd115_2 CB@21_mAd116_1 CB@21_mAd116_2 CB@21_mAd117_1 CB@21_mAd117_2 CB@21_mAd120_1 CB@21_mAd120_2 CB@21_mAd121_1 
+CB@21_mAd121_2 CB@21_mAd122_1 CB@21_mAd122_2 CB@21_mAd123_1 CB@21_mAd123_2 CB@21_mAd124_1 CB@21_mAd124_2 CB@21_mAd125_1 CB@21_mAd125_2 CB@21_mAd126_1 CB@21_mAd126_2 CB@21_mAd127_1 CB@21_mAd127_2 CB@21_mAd130_1 CB@21_mAd130_2 CB@21_mAd131_1 CB@21_mAd131_2 CB@21_mAd132_1 CB@21_mAd132_2 CB@21_mAd133_1 CB@21_mAd133_2 CB@21_mAd134_1 CB@21_mAd134_2 CB@21_mAd135_1 CB@21_mAd135_2 CB@21_mAd136_1 CB@21_mAd136_2 CB@21_mAd137_1 CB@21_mAd137_2 CB@21_mAd140_1 CB@21_mAd140_2 CB@21_mAd141_1 CB@21_mAd141_2 CB@21_mAd142_1 
+CB@21_mAd142_2 CB@21_mAd143_1 CB@21_mAd143_2 CB@21_mAd144_1 CB@21_mAd144_2 CB@21_mAd145_1 CB@21_mAd145_2 CB@21_mAd146_1 CB@21_mAd146_2 CB@21_mAd147_1 CB@21_mAd147_2 CB@21_mAd150_1 CB@21_mAd150_2 CB@21_mAd151_1 CB@21_mAd151_2 CB@21_mAd152_1 CB@21_mAd152_2 CB@21_mAd153_1 CB@21_mAd153_2 CB@21_mAd154_1 CB@21_mAd154_2 CB@21_mAd155_1 CB@21_mAd155_2 CB@21_mAd156_1 CB@21_mAd156_2 CB@21_mAd157_1 CB@21_mAd157_2 CB@21_mAd160_1 CB@21_mAd160_2 CB@21_mAd161_1 CB@21_mAd161_2 CB@21_mAd162_1 CB@21_mAd162_2 CB@21_mAd163_1 
+CB@21_mAd163_2 CB@21_mAd164_1 CB@21_mAd164_2 CB@21_mAd165_1 CB@21_mAd165_2 CB@21_mAd166_1 CB@21_mAd166_2 CB@21_mAd167_1 CB@21_mAd167_2 CB@21_mAd170_1 CB@21_mAd170_2 CB@21_mAd171_1 CB@21_mAd171_2 CB@21_mAd172_1 CB@21_mAd172_2 CB@21_mAd173_1 CB@21_mAd173_2 CB@21_mAd175_1 CB@21_mAd175_2 CB@21_mAd176_1 CB@21_mAd176_2 CB@21_mAd177_1 CB@21_mAd177_2 CB@21_mAd200_1 CB@21_mAd200_2 CB@21_mAd201_1 CB@21_mAd201_2 CB@21_mAd202_1 CB@21_mAd202_2 CB@21_mAd204_1 CB@21_mAd204_2 CB@21_mAd205_1 CB@21_mAd205_2 CB@21_mAd206_1 
+CB@21_mAd206_2 CB@21_mAd207_1 CB@21_mAd207_2 CB@21_mAd210_1 CB@21_mAd210_2 CB@21_mAd211_1 CB@21_mAd211_2 CB@21_mAd212_1 CB@21_mAd212_2 CB@21_mAd213_1 CB@21_mAd213_2 CB@21_mAd214_1 CB@21_mAd214_2 CB@21_mAd215_1 CB@21_mAd215_2 CB@21_mAd216_1 CB@21_mAd216_2 CB@21_mAd217_1 CB@21_mAd217_2 CB@21_mAd220_1 CB@21_mAd220_2 CB@21_mAd221_1 CB@21_mAd221_2 CB@21_mAd222_1 CB@21_mAd222_2 CB@21_mAd223_1 CB@21_mAd223_2 CB@21_mAd224_1 CB@21_mAd224_2 CB@21_mAd225_1 CB@21_mAd225_2 CB@21_mAd226_1 CB@21_mAd226_2 CB@21_mAd227_1 
+CB@21_mAd227_2 CB@21_mAd230_1 CB@21_mAd230_2 CB@21_mAd231_1 CB@21_mAd231_2 CB@21_mAd232_1 CB@21_mAd232_2 CB@21_mAd233_1 CB@21_mAd233_2 CB@21_mAd234_1 CB@21_mAd234_2 CB@21_mAd235_1 CB@21_mAd235_2 CB@21_mAd236_1 CB@21_mAd236_2 CB@21_mAd237_1 CB@21_mAd237_2 CB@21_mAd240_1 CB@21_mAd240_2 CB@21_mAd241_1 CB@21_mAd241_2 CB@21_mAd242_1 CB@21_mAd242_2 CB@21_mAd243_1 CB@21_mAd243_2 CB@21_mAd244_1 CB@21_mAd244_2 CB@21_mAd245_1 CB@21_mAd245_2 CB@21_mAd246_1 CB@21_mAd246_2 CB@21_mAd247_1 CB@21_mAd247_2 CB@21_mAd250_1 
+CB@21_mAd250_2 CB@21_mAd251_1 CB@21_mAd251_2 CB@21_mAd252_1 CB@21_mAd252_2 CB@21_mAd253_1 CB@21_mAd253_2 CB@21_mAd254_1 CB@21_mAd254_2 CB@21_mAd255_1 CB@21_mAd255_2 CB@21_mAd256_1 CB@21_mAd256_2 CB@21_mAd257_1 CB@21_mAd257_2 CB@21_mAd260_1 CB@21_mAd260_2 CB@21_mAd261_1 CB@21_mAd261_2 CB@21_mAd262_1 CB@21_mAd262_2 CB@21_mAd263_1 CB@21_mAd263_2 CB@21_mAd264_1 CB@21_mAd264_2 CB@21_mAd265_1 CB@21_mAd265_2 CB@21_mAd266_1 CB@21_mAd266_2 CB@21_mAd267_1 CB@21_mAd267_2 CB@21_mAd275_1 CB@21_mAd275_2 CB@21_mAd276_1 
+CB@21_mAd276_2 CB@21_mAd277_1 CB@21_mAd277_2 CB@21_mAd300_1 CB@21_mAd300_2 CB@21_mAd310_1 CB@21_mAd310_2 CB@21_mAd311_1 CB@21_mAd311_2 CB@21_mAd317_1 CB@21_mAd317_2 CB@21_mAd320_1 CB@21_mAd320_2 CB@21_mAd321_1 CB@21_mAd321_2 CB@21_mAd322_1 CB@21_mAd322_2 CB@21_mAd323_1 CB@21_mAd323_2 CB@21_mAd324_1 CB@21_mAd324_2 CB@21_mAd325_1 CB@21_mAd325_2 CB@21_mAd326_1 CB@21_mAd326_2 CB@21_mAd327_1 CB@21_mAd327_2 CB@21_mAd330_1 CB@21_mAd330_2 CB@21_mAd331_1 CB@21_mAd331_2 CB@21_mAd332_1 CB@21_mAd332_2 CB@21_mAd333_1 
+CB@21_mAd333_2 CB@21_mAd334_1 CB@21_mAd334_2 CB@21_mAd335_1 CB@21_mAd335_2 CB@21_mAd336_1 CB@21_mAd336_2 CB@21_mAd337_1 CB@21_mAd337_2 CB@21_mAd340_1 CB@21_mAd340_2 CB@21_mAd341_1 CB@21_mAd341_2 CB@21_mAd342_1 CB@21_mAd342_2 CB@21_mAd343_1 CB@21_mAd343_2 CB@21_mAd344_1 CB@21_mAd344_2 CB@21_mAd345_1 CB@21_mAd345_2 CB@21_mAd346_1 CB@21_mAd346_2 CB@21_mAd347_1 CB@21_mAd347_2 CB@21_mAd350_1 CB@21_mAd350_2 CB@21_mAd351_1 CB@21_mAd351_2 CB@21_mAd352_1 CB@21_mAd352_2 CB@21_mAd353_1 CB@21_mAd353_2 CB@21_mAd354_1 
+CB@21_mAd354_2 CB@21_mAd355_1 CB@21_mAd355_2 CB@21_mAd356_1 CB@21_mAd356_2 CB@21_mAd357_1 CB@21_mAd357_2 CB@21_mAd360_1 CB@21_mAd360_2 CB@21_mAd361_1 CB@21_mAd361_2 CB@21_mAd362_1 CB@21_mAd362_2 CB@21_mAd363_1 CB@21_mAd363_2 CB@21_mAd364_1 CB@21_mAd364_2 CB@21_mAd365_1 CB@21_mAd365_2 CB@21_mAd366_1 CB@21_mAd366_2 CB@21_mAd367_1 CB@21_mAd367_2 CB@21_mAd371_1 CB@21_mAd371_2 CB@21_mAd372_1 CB@21_mAd372_2 CB@21_mAd373_1 CB@21_mAd373_2 CB@21_mAd374_1 CB@21_mAd374_2 CB@21_mAd375_1 CB@21_mAd375_2 CB@21_mAd376_1 
+CB@21_mAd376_2 CB@21_mAd377_1 CB@21_mAd377_2 CB@21_mAd400_1 CB@21_mAd400_2 CB@21_mAd401_1 CB@21_mAd401_2 CB@21_mAd402_1 CB@21_mAd402_2 CB@21_mAd403_1 CB@21_mAd403_2 CB@21_mAd404_1 CB@21_mAd404_2 CB@21_mAd405_1 CB@21_mAd405_2 CB@21_mAd406_1 CB@21_mAd406_2 CB@21_mAd407_1 CB@21_mAd407_2 CB@21_mAd410_1 CB@21_mAd410_2 CB@21_mAd411_1 CB@21_mAd411_2 CB@21_mAd412_1 CB@21_mAd412_2 CB@21_mAd413_1 CB@21_mAd413_2 CB@21_mAd414_1 CB@21_mAd414_2 CB@21_mAd415_1 CB@21_mAd415_2 CB@21_mAd416_1 CB@21_mAd416_2 CB@21_mAd417_1 
+CB@21_mAd417_2 CB@21_mAd420_1 CB@21_mAd420_2 CB@21_mAd421_1 CB@21_mAd421_2 CB@21_mAd422_1 CB@21_mAd422_2 CB@21_mAd423_1 CB@21_mAd423_2 CB@21_mAd424_1 CB@21_mAd424_2 CB@21_mAd425_1 CB@21_mAd425_2 CB@21_mAd426_1 CB@21_mAd426_2 CB@21_mAd427_1 CB@21_mAd427_2 CB@21_mAd430_1 CB@21_mAd430_2 CB@21_mAd431_1 CB@21_mAd431_2 CB@21_mAd432_1 CB@21_mAd432_2 CB@21_mAd433_1 CB@21_mAd433_2 CB@21_mAd434_1 CB@21_mAd434_2 CB@21_mAd435_1 CB@21_mAd435_2 CB@21_mAd436_1 CB@21_mAd436_2 CB@21_mAd437_1 CB@21_mAd437_2 CB@21_mAd440_1 
+CB@21_mAd440_2 CB@21_mAd441_1 CB@21_mAd441_2 CB@21_mAd442_1 CB@21_mAd442_2 CB@21_mAd443_1 CB@21_mAd443_2 CB@21_mAd444_1 CB@21_mAd444_2 CB@21_mAd445_1 CB@21_mAd445_2 CB@21_mAd446_1 CB@21_mAd446_2 CB@21_mAd447_1 CB@21_mAd447_2 CB@21_mAd450_1 CB@21_mAd450_2 CB@21_mAd451_1 CB@21_mAd451_2 CB@21_mAd452_1 CB@21_mAd452_2 CB@21_mAd453_1 CB@21_mAd453_2 CB@21_mAd454_1 CB@21_mAd454_2 CB@21_mAd455_1 CB@21_mAd455_2 CB@21_mAd456_1 CB@21_mAd456_2 CB@21_mAd457_1 CB@21_mAd457_2 CB@21_mAd460_1 CB@21_mAd460_2 CB@21_mAd466_1 
+CB@21_mAd466_2 CB@21_mAd467_1 CB@21_mAd467_2 CB@21_mAd500_1 CB@21_mAd500_2 CB@21_mAd501_1 CB@21_mAd501_2 CB@21_mAd502_1 CB@21_mAd502_2 CB@21_mAd508_1 CB@21_mAd508_2 CB@21_mAd509_1 CB@21_mAd509_2 CB@21_mAd512_1 CB@21_mAd512_2 CB@21_mAd513_1 CB@21_mAd513_2 CB@21_mAd514_1 CB@21_mAd514_2 CB@21_mAd515_1 CB@21_mAd515_2 CB@21_mAd516_1 CB@21_mAd516_2 CB@21_mAd517_1 CB@21_mAd517_2 CB@21_mAd520_1 CB@21_mAd520_2 CB@21_mAd521_1 CB@21_mAd521_2 CB@21_mAd522_1 CB@21_mAd522_2 CB@21_mAd523_1 CB@21_mAd523_2 CB@21_mAd524_1 
+CB@21_mAd524_2 CB@21_mAd525_1 CB@21_mAd525_2 CB@21_mAd526_1 CB@21_mAd526_2 CB@21_mAd527_1 CB@21_mAd527_2 CB@21_mAd530_1 CB@21_mAd530_2 CB@21_mAd531_1 CB@21_mAd531_2 CB@21_mAd532_1 CB@21_mAd532_2 CB@21_mAd533_1 CB@21_mAd533_2 CB@21_mAd534_1 CB@21_mAd534_2 CB@21_mAd535_1 CB@21_mAd535_2 CB@21_mAd536_1 CB@21_mAd536_2 CB@21_mAd537_1 CB@21_mAd537_2 CB@21_mAd540_1 CB@21_mAd540_2 CB@21_mAd541_1 CB@21_mAd541_2 CB@21_mAd542_1 CB@21_mAd542_2 CB@21_mAd543_1 CB@21_mAd543_2 CB@21_mAd544_1 CB@21_mAd544_2 CB@21_mAd545_1 
+CB@21_mAd545_2 CB@21_mAd546_1 CB@21_mAd546_2 CB@21_mAd547_1 CB@21_mAd547_2 CB@21_mAd550_1 CB@21_mAd550_2 CB@21_mAd551_1 CB@21_mAd551_2 CB@21_mAd552_1 CB@21_mAd552_2 CB@21_mAd553_1 CB@21_mAd553_2 CB@21_mAd554_1 CB@21_mAd554_2 CB@21_mAd555_1 CB@21_mAd555_2 CB@21_mAd556_1 CB@21_mAd556_2 CB@21_mAd557_1 CB@21_mAd557_2 CB@21_mAd560_1 CB@21_mAd560_2 CB@21_mAd561_1 CB@21_mAd561_2 CB@21_mAd562_1 CB@21_mAd562_2 CB@21_mAd563_1 CB@21_mAd563_2 CB@21_mAd564_1 CB@21_mAd564_2 CB@21_mAd565_1 CB@21_mAd565_2 CB@21_mAd566_1 
+CB@21_mAd566_2 CB@21_mAd567_1 CB@21_mAd567_2 CB@21_mAd570_1 CB@21_mAd570_2 CB@21_mAd571_1 CB@21_mAd571_2 CB@21_mAd572_1 CB@21_mAd572_2 CB@21_mAd573_1 CB@21_mAd573_2 CB@21_mAd575_1 CB@21_mAd575_2 CB@21_mAd576_1 CB@21_mAd576_2 CB@21_mAd577_1 CB@21_mAd577_2 CB@21_mAd600_1 CB@21_mAd600_2 CB@21_mAd601_1 CB@21_mAd601_2 CB@21_mAd602_1 CB@21_mAd602_2 CB@21_mAd604_1 CB@21_mAd604_2 CB@21_mAd605_1 CB@21_mAd605_2 CB@21_mAd606_1 CB@21_mAd606_2 CB@21_mAd607_1 CB@21_mAd607_2 CB@21_mAd610_1 CB@21_mAd610_2 CB@21_mAd611_1 
+CB@21_mAd611_2 CB@21_mAd612_1 CB@21_mAd612_2 CB@21_mAd613_1 CB@21_mAd613_2 CB@21_mAd614_1 CB@21_mAd614_2 CB@21_mAd615_1 CB@21_mAd615_2 CB@21_mAd616_1 CB@21_mAd616_2 CB@21_mAd617_1 CB@21_mAd617_2 CB@21_mAd620_1 CB@21_mAd620_2 CB@21_mAd621_1 CB@21_mAd621_2 CB@21_mAd622_1 CB@21_mAd622_2 CB@21_mAd623_1 CB@21_mAd623_2 CB@21_mAd624_1 CB@21_mAd624_2 CB@21_mAd625_1 CB@21_mAd625_2 CB@21_mAd626_1 CB@21_mAd626_2 CB@21_mAd627_1 CB@21_mAd627_2 CB@21_mAd630_1 CB@21_mAd630_2 CB@21_mAd631_1 CB@21_mAd631_2 CB@21_mAd632_1 
+CB@21_mAd632_2 CB@21_mAd633_1 CB@21_mAd633_2 CB@21_mAd634_1 CB@21_mAd634_2 CB@21_mAd635_1 CB@21_mAd635_2 CB@21_mAd636_1 CB@21_mAd636_2 CB@21_mAd637_1 CB@21_mAd637_2 CB@21_mAd640_1 CB@21_mAd640_2 CB@21_mAd641_1 CB@21_mAd641_2 CB@21_mAd642_1 CB@21_mAd642_2 CB@21_mAd643_1 CB@21_mAd643_2 CB@21_mAd644_1 CB@21_mAd644_2 CB@21_mAd645_1 CB@21_mAd645_2 CB@21_mAd646_1 CB@21_mAd646_2 CB@21_mAd647_1 CB@21_mAd647_2 CB@21_mAd650_1 CB@21_mAd650_2 CB@21_mAd651_1 CB@21_mAd651_2 CB@21_mAd652_1 CB@21_mAd652_2 CB@21_mAd653_1 
+CB@21_mAd653_2 CB@21_mAd654_1 CB@21_mAd654_2 CB@21_mAd655_1 CB@21_mAd655_2 CB@21_mAd656_1 CB@21_mAd656_2 CB@21_mAd657_1 CB@21_mAd657_2 CB@21_mAd660_1 CB@21_mAd660_2 CB@21_mAd661_1 CB@21_mAd661_2 CB@21_mAd662_1 CB@21_mAd662_2 CB@21_mAd663_1 CB@21_mAd663_2 CB@21_mAd664_1 CB@21_mAd664_2 CB@21_mAd665_1 CB@21_mAd665_2 CB@21_mAd666_1 CB@21_mAd666_2 CB@21_mAd667_1 CB@21_mAd667_2 CB@21_mAd675_1 CB@21_mAd675_2 CB@21_mAd676_1 CB@21_mAd676_2 CB@21_mAd677_1 CB@21_mAd677_2 CB@21_mAd700_1 CB@21_mAd700_2 CB@21_mAd710_1 
+CB@21_mAd710_2 CB@21_mAd711_1 CB@21_mAd711_2 CB@21_mAd717_1 CB@21_mAd717_2 CB@21_mAd720_1 CB@21_mAd720_2 CB@21_mAd721_1 CB@21_mAd721_2 CB@21_mAd722_1 CB@21_mAd722_2 CB@21_mAd723_1 CB@21_mAd723_2 CB@21_mAd724_1 CB@21_mAd724_2 CB@21_mAd725_1 CB@21_mAd725_2 CB@21_mAd726_1 CB@21_mAd726_2 CB@21_mAd727_1 CB@21_mAd727_2 CB@21_mAd730_1 CB@21_mAd730_2 CB@21_mAd731_1 CB@21_mAd731_2 CB@21_mAd732_1 CB@21_mAd732_2 CB@21_mAd733_1 CB@21_mAd733_2 CB@21_mAd734_1 CB@21_mAd734_2 CB@21_mAd735_1 CB@21_mAd735_2 CB@21_mAd736_1 
+CB@21_mAd736_2 CB@21_mAd737_1 CB@21_mAd737_2 CB@21_mAd740_1 CB@21_mAd740_2 CB@21_mAd741_1 CB@21_mAd741_2 CB@21_mAd742_1 CB@21_mAd742_2 CB@21_mAd743_1 CB@21_mAd743_2 CB@21_mAd744_1 CB@21_mAd744_2 CB@21_mAd745_1 CB@21_mAd745_2 CB@21_mAd746_1 CB@21_mAd746_2 CB@21_mAd747_1 CB@21_mAd747_2 CB@21_mAd750_1 CB@21_mAd750_2 CB@21_mAd751_1 CB@21_mAd751_2 CB@21_mAd752_1 CB@21_mAd752_2 CB@21_mAd753_1 CB@21_mAd753_2 CB@21_mAd754_1 CB@21_mAd754_2 CB@21_mAd755_1 CB@21_mAd755_2 CB@21_mAd756_1 CB@21_mAd756_2 CB@21_mAd757_1 
+CB@21_mAd757_2 CB@21_mAd760_1 CB@21_mAd760_2 CB@21_mAd761_1 CB@21_mAd761_2 CB@21_mAd762_1 CB@21_mAd762_2 CB@21_mAd763_1 CB@21_mAd763_2 CB@21_mAd764_1 CB@21_mAd764_2 CB@21_mAd765_1 CB@21_mAd765_2 CB@21_mAd766_1 CB@21_mAd766_2 CB@21_mAd767_1 CB@21_mAd767_2 CB@21_mAd771_1 CB@21_mAd771_2 CB@21_mAd772_1 CB@21_mAd772_2 CB@21_mAd773_1 CB@21_mAd773_2 CB@21_mAd774_1 CB@21_mAd774_2 CB@21_mAd775_1 CB@21_mAd775_2 CB@21_mAd776_1 CB@21_mAd776_2 CB@21_mAd777_1 CB@21_mAd777_2 CB@21_X0 CB@21_X1 CB@21_X10 CB@21_X11 
+CB@21_X12 CB@21_X13 CB@21_X2 CB@21_X3 CB@21_X4 CB@21_X5 CB@21_X6 CB@21_X7 CB@21_X8 CB@21_X9 CB@21_Y1 CB@21_Y10 CB@21_Y11 CB@21_Y12 CB@21_Y2 CB@21_Y3 CB@21_Y4 CB@21_Y5 CB@21_Y6 CB@21_Y7 CB@21_Y8 CB@21_Y9 CB@21_Z1 CB@21_Z10 CB@21_Z11 CB@21_Z12 CB@21_Z2 CB@21_Z3 CB@21_Z4 CB@21_Z5 CB@21_Z6 CB@21_Z7 CB@21_Z8 CB@21_Z9 _5400TP094__CB
XCB@22 CB@22_K0 CB@22_K1 CB@22_K10 CB@22_K11 CB@22_K12 CB@22_K13 CB@22_K2 CB@22_K3 CB@22_K4 CB@22_K5 CB@22_K6 CB@22_K7 CB@22_K8 CB@22_K9 CB@22_mAd000_1 CB@22_mAd000_2 CB@22_mAd001_1 CB@22_mAd001_2 CB@22_mAd002_1 CB@22_mAd002_2 CB@22_mAd003_1 CB@22_mAd003_2 CB@22_mAd004_1 CB@22_mAd004_2 CB@22_mAd005_1 CB@22_mAd005_2 CB@22_mAd006_1 CB@22_mAd006_2 CB@22_mAd007_1 CB@22_mAd007_2 CB@22_mAd010_1 CB@22_mAd010_2 CB@22_mAd011_1 CB@22_mAd011_2 CB@22_mAd012_1 CB@22_mAd012_2 CB@22_mAd013_1 CB@22_mAd013_2 CB@22_mAd014_1 
+CB@22_mAd014_2 CB@22_mAd015_1 CB@22_mAd015_2 CB@22_mAd016_1 CB@22_mAd016_2 CB@22_mAd017_1 CB@22_mAd017_2 CB@22_mAd020_1 CB@22_mAd020_2 CB@22_mAd021_1 CB@22_mAd021_2 CB@22_mAd022_1 CB@22_mAd022_2 CB@22_mAd023_1 CB@22_mAd023_2 CB@22_mAd024_1 CB@22_mAd024_2 CB@22_mAd025_1 CB@22_mAd025_2 CB@22_mAd026_1 CB@22_mAd026_2 CB@22_mAd027_1 CB@22_mAd027_2 CB@22_mAd030_1 CB@22_mAd030_2 CB@22_mAd031_1 CB@22_mAd031_2 CB@22_mAd032_1 CB@22_mAd032_2 CB@22_mAd033_1 CB@22_mAd033_2 CB@22_mAd034_1 CB@22_mAd034_2 CB@22_mAd035_1 
+CB@22_mAd035_2 CB@22_mAd036_1 CB@22_mAd036_2 CB@22_mAd037_1 CB@22_mAd037_2 CB@22_mAd040_1 CB@22_mAd040_2 CB@22_mAd041_1 CB@22_mAd041_2 CB@22_mAd042_1 CB@22_mAd042_2 CB@22_mAd043_1 CB@22_mAd043_2 CB@22_mAd044_1 CB@22_mAd044_2 CB@22_mAd045_1 CB@22_mAd045_2 CB@22_mAd046_1 CB@22_mAd046_2 CB@22_mAd047_1 CB@22_mAd047_2 CB@22_mAd050_1 CB@22_mAd050_2 CB@22_mAd051_1 CB@22_mAd051_2 CB@22_mAd052_1 CB@22_mAd052_2 CB@22_mAd053_1 CB@22_mAd053_2 CB@22_mAd054_1 CB@22_mAd054_2 CB@22_mAd055_1 CB@22_mAd055_2 CB@22_mAd056_1 
+CB@22_mAd056_2 CB@22_mAd057_1 CB@22_mAd057_2 CB@22_mAd060_1 CB@22_mAd060_2 CB@22_mAd066_1 CB@22_mAd066_2 CB@22_mAd067_1 CB@22_mAd067_2 CB@22_mAd100_1 CB@22_mAd100_2 CB@22_mAd101_1 CB@22_mAd101_2 CB@22_mAd102_1 CB@22_mAd102_2 CB@22_mAd110_1 CB@22_mAd110_2 CB@22_mAd111_1 CB@22_mAd111_2 CB@22_mAd112_1 CB@22_mAd112_2 CB@22_mAd113_1 CB@22_mAd113_2 CB@22_mAd114_1 CB@22_mAd114_2 CB@22_mAd115_1 CB@22_mAd115_2 CB@22_mAd116_1 CB@22_mAd116_2 CB@22_mAd117_1 CB@22_mAd117_2 CB@22_mAd120_1 CB@22_mAd120_2 CB@22_mAd121_1 
+CB@22_mAd121_2 CB@22_mAd122_1 CB@22_mAd122_2 CB@22_mAd123_1 CB@22_mAd123_2 CB@22_mAd124_1 CB@22_mAd124_2 CB@22_mAd125_1 CB@22_mAd125_2 CB@22_mAd126_1 CB@22_mAd126_2 CB@22_mAd127_1 CB@22_mAd127_2 CB@22_mAd130_1 CB@22_mAd130_2 CB@22_mAd131_1 CB@22_mAd131_2 CB@22_mAd132_1 CB@22_mAd132_2 CB@22_mAd133_1 CB@22_mAd133_2 CB@22_mAd134_1 CB@22_mAd134_2 CB@22_mAd135_1 CB@22_mAd135_2 CB@22_mAd136_1 CB@22_mAd136_2 CB@22_mAd137_1 CB@22_mAd137_2 CB@22_mAd140_1 CB@22_mAd140_2 CB@22_mAd141_1 CB@22_mAd141_2 CB@22_mAd142_1 
+CB@22_mAd142_2 CB@22_mAd143_1 CB@22_mAd143_2 CB@22_mAd144_1 CB@22_mAd144_2 CB@22_mAd145_1 CB@22_mAd145_2 CB@22_mAd146_1 CB@22_mAd146_2 CB@22_mAd147_1 CB@22_mAd147_2 CB@22_mAd150_1 CB@22_mAd150_2 CB@22_mAd151_1 CB@22_mAd151_2 CB@22_mAd152_1 CB@22_mAd152_2 CB@22_mAd153_1 CB@22_mAd153_2 CB@22_mAd154_1 CB@22_mAd154_2 CB@22_mAd155_1 CB@22_mAd155_2 CB@22_mAd156_1 CB@22_mAd156_2 CB@22_mAd157_1 CB@22_mAd157_2 CB@22_mAd160_1 CB@22_mAd160_2 CB@22_mAd161_1 CB@22_mAd161_2 CB@22_mAd162_1 CB@22_mAd162_2 CB@22_mAd163_1 
+CB@22_mAd163_2 CB@22_mAd164_1 CB@22_mAd164_2 CB@22_mAd165_1 CB@22_mAd165_2 CB@22_mAd166_1 CB@22_mAd166_2 CB@22_mAd167_1 CB@22_mAd167_2 CB@22_mAd170_1 CB@22_mAd170_2 CB@22_mAd171_1 CB@22_mAd171_2 CB@22_mAd172_1 CB@22_mAd172_2 CB@22_mAd173_1 CB@22_mAd173_2 CB@22_mAd175_1 CB@22_mAd175_2 CB@22_mAd176_1 CB@22_mAd176_2 CB@22_mAd177_1 CB@22_mAd177_2 CB@22_mAd200_1 CB@22_mAd200_2 CB@22_mAd201_1 CB@22_mAd201_2 CB@22_mAd202_1 CB@22_mAd202_2 CB@22_mAd204_1 CB@22_mAd204_2 CB@22_mAd205_1 CB@22_mAd205_2 CB@22_mAd206_1 
+CB@22_mAd206_2 CB@22_mAd207_1 CB@22_mAd207_2 CB@22_mAd210_1 CB@22_mAd210_2 CB@22_mAd211_1 CB@22_mAd211_2 CB@22_mAd212_1 CB@22_mAd212_2 CB@22_mAd213_1 CB@22_mAd213_2 CB@22_mAd214_1 CB@22_mAd214_2 CB@22_mAd215_1 CB@22_mAd215_2 CB@22_mAd216_1 CB@22_mAd216_2 CB@22_mAd217_1 CB@22_mAd217_2 CB@22_mAd220_1 CB@22_mAd220_2 CB@22_mAd221_1 CB@22_mAd221_2 CB@22_mAd222_1 CB@22_mAd222_2 CB@22_mAd223_1 CB@22_mAd223_2 CB@22_mAd224_1 CB@22_mAd224_2 CB@22_mAd225_1 CB@22_mAd225_2 CB@22_mAd226_1 CB@22_mAd226_2 CB@22_mAd227_1 
+CB@22_mAd227_2 CB@22_mAd230_1 CB@22_mAd230_2 CB@22_mAd231_1 CB@22_mAd231_2 CB@22_mAd232_1 CB@22_mAd232_2 CB@22_mAd233_1 CB@22_mAd233_2 CB@22_mAd234_1 CB@22_mAd234_2 CB@22_mAd235_1 CB@22_mAd235_2 CB@22_mAd236_1 CB@22_mAd236_2 CB@22_mAd237_1 CB@22_mAd237_2 CB@22_mAd240_1 CB@22_mAd240_2 CB@22_mAd241_1 CB@22_mAd241_2 CB@22_mAd242_1 CB@22_mAd242_2 CB@22_mAd243_1 CB@22_mAd243_2 CB@22_mAd244_1 CB@22_mAd244_2 CB@22_mAd245_1 CB@22_mAd245_2 CB@22_mAd246_1 CB@22_mAd246_2 CB@22_mAd247_1 CB@22_mAd247_2 CB@22_mAd250_1 
+CB@22_mAd250_2 CB@22_mAd251_1 CB@22_mAd251_2 CB@22_mAd252_1 CB@22_mAd252_2 CB@22_mAd253_1 CB@22_mAd253_2 CB@22_mAd254_1 CB@22_mAd254_2 CB@22_mAd255_1 CB@22_mAd255_2 CB@22_mAd256_1 CB@22_mAd256_2 CB@22_mAd257_1 CB@22_mAd257_2 CB@22_mAd260_1 CB@22_mAd260_2 CB@22_mAd261_1 CB@22_mAd261_2 CB@22_mAd262_1 CB@22_mAd262_2 CB@22_mAd263_1 CB@22_mAd263_2 CB@22_mAd264_1 CB@22_mAd264_2 CB@22_mAd265_1 CB@22_mAd265_2 CB@22_mAd266_1 CB@22_mAd266_2 CB@22_mAd267_1 CB@22_mAd267_2 CB@22_mAd275_1 CB@22_mAd275_2 CB@22_mAd276_1 
+CB@22_mAd276_2 CB@22_mAd277_1 CB@22_mAd277_2 CB@22_mAd300_1 CB@22_mAd300_2 CB@22_mAd310_1 CB@22_mAd310_2 CB@22_mAd311_1 CB@22_mAd311_2 CB@22_mAd317_1 CB@22_mAd317_2 CB@22_mAd320_1 CB@22_mAd320_2 CB@22_mAd321_1 CB@22_mAd321_2 CB@22_mAd322_1 CB@22_mAd322_2 CB@22_mAd323_1 CB@22_mAd323_2 CB@22_mAd324_1 CB@22_mAd324_2 CB@22_mAd325_1 CB@22_mAd325_2 CB@22_mAd326_1 CB@22_mAd326_2 CB@22_mAd327_1 CB@22_mAd327_2 CB@22_mAd330_1 CB@22_mAd330_2 CB@22_mAd331_1 CB@22_mAd331_2 CB@22_mAd332_1 CB@22_mAd332_2 CB@22_mAd333_1 
+CB@22_mAd333_2 CB@22_mAd334_1 CB@22_mAd334_2 CB@22_mAd335_1 CB@22_mAd335_2 CB@22_mAd336_1 CB@22_mAd336_2 CB@22_mAd337_1 CB@22_mAd337_2 CB@22_mAd340_1 CB@22_mAd340_2 CB@22_mAd341_1 CB@22_mAd341_2 CB@22_mAd342_1 CB@22_mAd342_2 CB@22_mAd343_1 CB@22_mAd343_2 CB@22_mAd344_1 CB@22_mAd344_2 CB@22_mAd345_1 CB@22_mAd345_2 CB@22_mAd346_1 CB@22_mAd346_2 CB@22_mAd347_1 CB@22_mAd347_2 CB@22_mAd350_1 CB@22_mAd350_2 CB@22_mAd351_1 CB@22_mAd351_2 CB@22_mAd352_1 CB@22_mAd352_2 CB@22_mAd353_1 CB@22_mAd353_2 CB@22_mAd354_1 
+CB@22_mAd354_2 CB@22_mAd355_1 CB@22_mAd355_2 CB@22_mAd356_1 CB@22_mAd356_2 CB@22_mAd357_1 CB@22_mAd357_2 CB@22_mAd360_1 CB@22_mAd360_2 CB@22_mAd361_1 CB@22_mAd361_2 CB@22_mAd362_1 CB@22_mAd362_2 CB@22_mAd363_1 CB@22_mAd363_2 CB@22_mAd364_1 CB@22_mAd364_2 CB@22_mAd365_1 CB@22_mAd365_2 CB@22_mAd366_1 CB@22_mAd366_2 CB@22_mAd367_1 CB@22_mAd367_2 CB@22_mAd371_1 CB@22_mAd371_2 CB@22_mAd372_1 CB@22_mAd372_2 CB@22_mAd373_1 CB@22_mAd373_2 CB@22_mAd374_1 CB@22_mAd374_2 CB@22_mAd375_1 CB@22_mAd375_2 CB@22_mAd376_1 
+CB@22_mAd376_2 CB@22_mAd377_1 CB@22_mAd377_2 CB@22_mAd400_1 CB@22_mAd400_2 CB@22_mAd401_1 CB@22_mAd401_2 CB@22_mAd402_1 CB@22_mAd402_2 CB@22_mAd403_1 CB@22_mAd403_2 CB@22_mAd404_1 CB@22_mAd404_2 CB@22_mAd405_1 CB@22_mAd405_2 CB@22_mAd406_1 CB@22_mAd406_2 CB@22_mAd407_1 CB@22_mAd407_2 CB@22_mAd410_1 CB@22_mAd410_2 CB@22_mAd411_1 CB@22_mAd411_2 CB@22_mAd412_1 CB@22_mAd412_2 CB@22_mAd413_1 CB@22_mAd413_2 CB@22_mAd414_1 CB@22_mAd414_2 CB@22_mAd415_1 CB@22_mAd415_2 CB@22_mAd416_1 CB@22_mAd416_2 CB@22_mAd417_1 
+CB@22_mAd417_2 CB@22_mAd420_1 CB@22_mAd420_2 CB@22_mAd421_1 CB@22_mAd421_2 CB@22_mAd422_1 CB@22_mAd422_2 CB@22_mAd423_1 CB@22_mAd423_2 CB@22_mAd424_1 CB@22_mAd424_2 CB@22_mAd425_1 CB@22_mAd425_2 CB@22_mAd426_1 CB@22_mAd426_2 CB@22_mAd427_1 CB@22_mAd427_2 CB@22_mAd430_1 CB@22_mAd430_2 CB@22_mAd431_1 CB@22_mAd431_2 CB@22_mAd432_1 CB@22_mAd432_2 CB@22_mAd433_1 CB@22_mAd433_2 CB@22_mAd434_1 CB@22_mAd434_2 CB@22_mAd435_1 CB@22_mAd435_2 CB@22_mAd436_1 CB@22_mAd436_2 CB@22_mAd437_1 CB@22_mAd437_2 CB@22_mAd440_1 
+CB@22_mAd440_2 CB@22_mAd441_1 CB@22_mAd441_2 CB@22_mAd442_1 CB@22_mAd442_2 CB@22_mAd443_1 CB@22_mAd443_2 CB@22_mAd444_1 CB@22_mAd444_2 CB@22_mAd445_1 CB@22_mAd445_2 CB@22_mAd446_1 CB@22_mAd446_2 CB@22_mAd447_1 CB@22_mAd447_2 CB@22_mAd450_1 CB@22_mAd450_2 CB@22_mAd451_1 CB@22_mAd451_2 CB@22_mAd452_1 CB@22_mAd452_2 CB@22_mAd453_1 CB@22_mAd453_2 CB@22_mAd454_1 CB@22_mAd454_2 CB@22_mAd455_1 CB@22_mAd455_2 CB@22_mAd456_1 CB@22_mAd456_2 CB@22_mAd457_1 CB@22_mAd457_2 CB@22_mAd460_1 CB@22_mAd460_2 CB@22_mAd466_1 
+CB@22_mAd466_2 CB@22_mAd467_1 CB@22_mAd467_2 CB@22_mAd500_1 CB@22_mAd500_2 CB@22_mAd501_1 CB@22_mAd501_2 CB@22_mAd502_1 CB@22_mAd502_2 CB@22_mAd508_1 CB@22_mAd508_2 CB@22_mAd509_1 CB@22_mAd509_2 CB@22_mAd512_1 CB@22_mAd512_2 CB@22_mAd513_1 CB@22_mAd513_2 CB@22_mAd514_1 CB@22_mAd514_2 CB@22_mAd515_1 CB@22_mAd515_2 CB@22_mAd516_1 CB@22_mAd516_2 CB@22_mAd517_1 CB@22_mAd517_2 CB@22_mAd520_1 CB@22_mAd520_2 CB@22_mAd521_1 CB@22_mAd521_2 CB@22_mAd522_1 CB@22_mAd522_2 CB@22_mAd523_1 CB@22_mAd523_2 CB@22_mAd524_1 
+CB@22_mAd524_2 CB@22_mAd525_1 CB@22_mAd525_2 CB@22_mAd526_1 CB@22_mAd526_2 CB@22_mAd527_1 CB@22_mAd527_2 CB@22_mAd530_1 CB@22_mAd530_2 CB@22_mAd531_1 CB@22_mAd531_2 CB@22_mAd532_1 CB@22_mAd532_2 CB@22_mAd533_1 CB@22_mAd533_2 CB@22_mAd534_1 CB@22_mAd534_2 CB@22_mAd535_1 CB@22_mAd535_2 CB@22_mAd536_1 CB@22_mAd536_2 CB@22_mAd537_1 CB@22_mAd537_2 CB@22_mAd540_1 CB@22_mAd540_2 CB@22_mAd541_1 CB@22_mAd541_2 CB@22_mAd542_1 CB@22_mAd542_2 CB@22_mAd543_1 CB@22_mAd543_2 CB@22_mAd544_1 CB@22_mAd544_2 CB@22_mAd545_1 
+CB@22_mAd545_2 CB@22_mAd546_1 CB@22_mAd546_2 CB@22_mAd547_1 CB@22_mAd547_2 CB@22_mAd550_1 CB@22_mAd550_2 CB@22_mAd551_1 CB@22_mAd551_2 CB@22_mAd552_1 CB@22_mAd552_2 CB@22_mAd553_1 CB@22_mAd553_2 CB@22_mAd554_1 CB@22_mAd554_2 CB@22_mAd555_1 CB@22_mAd555_2 CB@22_mAd556_1 CB@22_mAd556_2 CB@22_mAd557_1 CB@22_mAd557_2 CB@22_mAd560_1 CB@22_mAd560_2 CB@22_mAd561_1 CB@22_mAd561_2 CB@22_mAd562_1 CB@22_mAd562_2 CB@22_mAd563_1 CB@22_mAd563_2 CB@22_mAd564_1 CB@22_mAd564_2 CB@22_mAd565_1 CB@22_mAd565_2 CB@22_mAd566_1 
+CB@22_mAd566_2 CB@22_mAd567_1 CB@22_mAd567_2 CB@22_mAd570_1 CB@22_mAd570_2 CB@22_mAd571_1 CB@22_mAd571_2 CB@22_mAd572_1 CB@22_mAd572_2 CB@22_mAd573_1 CB@22_mAd573_2 CB@22_mAd575_1 CB@22_mAd575_2 CB@22_mAd576_1 CB@22_mAd576_2 CB@22_mAd577_1 CB@22_mAd577_2 CB@22_mAd600_1 CB@22_mAd600_2 CB@22_mAd601_1 CB@22_mAd601_2 CB@22_mAd602_1 CB@22_mAd602_2 CB@22_mAd604_1 CB@22_mAd604_2 CB@22_mAd605_1 CB@22_mAd605_2 CB@22_mAd606_1 CB@22_mAd606_2 CB@22_mAd607_1 CB@22_mAd607_2 CB@22_mAd610_1 CB@22_mAd610_2 CB@22_mAd611_1 
+CB@22_mAd611_2 CB@22_mAd612_1 CB@22_mAd612_2 CB@22_mAd613_1 CB@22_mAd613_2 CB@22_mAd614_1 CB@22_mAd614_2 CB@22_mAd615_1 CB@22_mAd615_2 CB@22_mAd616_1 CB@22_mAd616_2 CB@22_mAd617_1 CB@22_mAd617_2 CB@22_mAd620_1 CB@22_mAd620_2 CB@22_mAd621_1 CB@22_mAd621_2 CB@22_mAd622_1 CB@22_mAd622_2 CB@22_mAd623_1 CB@22_mAd623_2 CB@22_mAd624_1 CB@22_mAd624_2 CB@22_mAd625_1 CB@22_mAd625_2 CB@22_mAd626_1 CB@22_mAd626_2 CB@22_mAd627_1 CB@22_mAd627_2 CB@22_mAd630_1 CB@22_mAd630_2 CB@22_mAd631_1 CB@22_mAd631_2 CB@22_mAd632_1 
+CB@22_mAd632_2 CB@22_mAd633_1 CB@22_mAd633_2 CB@22_mAd634_1 CB@22_mAd634_2 CB@22_mAd635_1 CB@22_mAd635_2 CB@22_mAd636_1 CB@22_mAd636_2 CB@22_mAd637_1 CB@22_mAd637_2 CB@22_mAd640_1 CB@22_mAd640_2 CB@22_mAd641_1 CB@22_mAd641_2 CB@22_mAd642_1 CB@22_mAd642_2 CB@22_mAd643_1 CB@22_mAd643_2 CB@22_mAd644_1 CB@22_mAd644_2 CB@22_mAd645_1 CB@22_mAd645_2 CB@22_mAd646_1 CB@22_mAd646_2 CB@22_mAd647_1 CB@22_mAd647_2 CB@22_mAd650_1 CB@22_mAd650_2 CB@22_mAd651_1 CB@22_mAd651_2 CB@22_mAd652_1 CB@22_mAd652_2 CB@22_mAd653_1 
+CB@22_mAd653_2 CB@22_mAd654_1 CB@22_mAd654_2 CB@22_mAd655_1 CB@22_mAd655_2 CB@22_mAd656_1 CB@22_mAd656_2 CB@22_mAd657_1 CB@22_mAd657_2 CB@22_mAd660_1 CB@22_mAd660_2 CB@22_mAd661_1 CB@22_mAd661_2 CB@22_mAd662_1 CB@22_mAd662_2 CB@22_mAd663_1 CB@22_mAd663_2 CB@22_mAd664_1 CB@22_mAd664_2 CB@22_mAd665_1 CB@22_mAd665_2 CB@22_mAd666_1 CB@22_mAd666_2 CB@22_mAd667_1 CB@22_mAd667_2 CB@22_mAd675_1 CB@22_mAd675_2 CB@22_mAd676_1 CB@22_mAd676_2 CB@22_mAd677_1 CB@22_mAd677_2 CB@22_mAd700_1 CB@22_mAd700_2 CB@22_mAd710_1 
+CB@22_mAd710_2 CB@22_mAd711_1 CB@22_mAd711_2 CB@22_mAd717_1 CB@22_mAd717_2 CB@22_mAd720_1 CB@22_mAd720_2 CB@22_mAd721_1 CB@22_mAd721_2 CB@22_mAd722_1 CB@22_mAd722_2 CB@22_mAd723_1 CB@22_mAd723_2 CB@22_mAd724_1 CB@22_mAd724_2 CB@22_mAd725_1 CB@22_mAd725_2 CB@22_mAd726_1 CB@22_mAd726_2 CB@22_mAd727_1 CB@22_mAd727_2 CB@22_mAd730_1 CB@22_mAd730_2 CB@22_mAd731_1 CB@22_mAd731_2 CB@22_mAd732_1 CB@22_mAd732_2 CB@22_mAd733_1 CB@22_mAd733_2 CB@22_mAd734_1 CB@22_mAd734_2 CB@22_mAd735_1 CB@22_mAd735_2 CB@22_mAd736_1 
+CB@22_mAd736_2 CB@22_mAd737_1 CB@22_mAd737_2 CB@22_mAd740_1 CB@22_mAd740_2 CB@22_mAd741_1 CB@22_mAd741_2 CB@22_mAd742_1 CB@22_mAd742_2 CB@22_mAd743_1 CB@22_mAd743_2 CB@22_mAd744_1 CB@22_mAd744_2 CB@22_mAd745_1 CB@22_mAd745_2 CB@22_mAd746_1 CB@22_mAd746_2 CB@22_mAd747_1 CB@22_mAd747_2 CB@22_mAd750_1 CB@22_mAd750_2 CB@22_mAd751_1 CB@22_mAd751_2 CB@22_mAd752_1 CB@22_mAd752_2 CB@22_mAd753_1 CB@22_mAd753_2 CB@22_mAd754_1 CB@22_mAd754_2 CB@22_mAd755_1 CB@22_mAd755_2 CB@22_mAd756_1 CB@22_mAd756_2 CB@22_mAd757_1 
+CB@22_mAd757_2 CB@22_mAd760_1 CB@22_mAd760_2 CB@22_mAd761_1 CB@22_mAd761_2 CB@22_mAd762_1 CB@22_mAd762_2 CB@22_mAd763_1 CB@22_mAd763_2 CB@22_mAd764_1 CB@22_mAd764_2 CB@22_mAd765_1 CB@22_mAd765_2 CB@22_mAd766_1 CB@22_mAd766_2 CB@22_mAd767_1 CB@22_mAd767_2 CB@22_mAd771_1 CB@22_mAd771_2 CB@22_mAd772_1 CB@22_mAd772_2 CB@22_mAd773_1 CB@22_mAd773_2 CB@22_mAd774_1 CB@22_mAd774_2 CB@22_mAd775_1 CB@22_mAd775_2 CB@22_mAd776_1 CB@22_mAd776_2 CB@22_mAd777_1 CB@22_mAd777_2 CB@22_X0 CB@22_X1 CB@22_X10 CB@22_X11 
+CB@22_X12 CB@22_X13 CB@22_X2 CB@22_X3 CB@22_X4 CB@22_X5 CB@22_X6 CB@22_X7 CB@22_X8 CB@22_X9 CB@22_Y1 CB@22_Y10 CB@22_Y11 CB@22_Y12 CB@22_Y2 CB@22_Y3 CB@22_Y4 CB@22_Y5 CB@22_Y6 CB@22_Y7 CB@22_Y8 CB@22_Y9 CB@22_Z1 CB@22_Z10 CB@22_Z11 CB@22_Z12 CB@22_Z2 CB@22_Z3 CB@22_Z4 CB@22_Z5 CB@22_Z6 CB@22_Z7 CB@22_Z8 CB@22_Z9 _5400TP094__CB
XCB@23 CB@23_K0 CB@23_K1 CB@23_K10 CB@23_K11 CB@23_K12 CB@23_K13 CB@23_K2 CB@23_K3 CB@23_K4 CB@23_K5 CB@23_K6 CB@23_K7 CB@23_K8 CB@23_K9 CB@23_mAd000_1 CB@23_mAd000_2 CB@23_mAd001_1 CB@23_mAd001_2 CB@23_mAd002_1 CB@23_mAd002_2 CB@23_mAd003_1 CB@23_mAd003_2 CB@23_mAd004_1 CB@23_mAd004_2 CB@23_mAd005_1 CB@23_mAd005_2 CB@23_mAd006_1 CB@23_mAd006_2 CB@23_mAd007_1 CB@23_mAd007_2 CB@23_mAd010_1 CB@23_mAd010_2 CB@23_mAd011_1 CB@23_mAd011_2 CB@23_mAd012_1 CB@23_mAd012_2 CB@23_mAd013_1 CB@23_mAd013_2 CB@23_mAd014_1 
+CB@23_mAd014_2 CB@23_mAd015_1 CB@23_mAd015_2 CB@23_mAd016_1 CB@23_mAd016_2 CB@23_mAd017_1 CB@23_mAd017_2 CB@23_mAd020_1 CB@23_mAd020_2 CB@23_mAd021_1 CB@23_mAd021_2 CB@23_mAd022_1 CB@23_mAd022_2 CB@23_mAd023_1 CB@23_mAd023_2 CB@23_mAd024_1 CB@23_mAd024_2 CB@23_mAd025_1 CB@23_mAd025_2 CB@23_mAd026_1 CB@23_mAd026_2 CB@23_mAd027_1 CB@23_mAd027_2 CB@23_mAd030_1 CB@23_mAd030_2 CB@23_mAd031_1 CB@23_mAd031_2 CB@23_mAd032_1 CB@23_mAd032_2 CB@23_mAd033_1 CB@23_mAd033_2 CB@23_mAd034_1 CB@23_mAd034_2 CB@23_mAd035_1 
+CB@23_mAd035_2 CB@23_mAd036_1 CB@23_mAd036_2 CB@23_mAd037_1 CB@23_mAd037_2 CB@23_mAd040_1 CB@23_mAd040_2 CB@23_mAd041_1 CB@23_mAd041_2 CB@23_mAd042_1 CB@23_mAd042_2 CB@23_mAd043_1 CB@23_mAd043_2 CB@23_mAd044_1 CB@23_mAd044_2 CB@23_mAd045_1 CB@23_mAd045_2 CB@23_mAd046_1 CB@23_mAd046_2 CB@23_mAd047_1 CB@23_mAd047_2 CB@23_mAd050_1 CB@23_mAd050_2 CB@23_mAd051_1 CB@23_mAd051_2 CB@23_mAd052_1 CB@23_mAd052_2 CB@23_mAd053_1 CB@23_mAd053_2 CB@23_mAd054_1 CB@23_mAd054_2 CB@23_mAd055_1 CB@23_mAd055_2 CB@23_mAd056_1 
+CB@23_mAd056_2 CB@23_mAd057_1 CB@23_mAd057_2 CB@23_mAd060_1 CB@23_mAd060_2 CB@23_mAd066_1 CB@23_mAd066_2 CB@23_mAd067_1 CB@23_mAd067_2 CB@23_mAd100_1 CB@23_mAd100_2 CB@23_mAd101_1 CB@23_mAd101_2 CB@23_mAd102_1 CB@23_mAd102_2 CB@23_mAd110_1 CB@23_mAd110_2 CB@23_mAd111_1 CB@23_mAd111_2 CB@23_mAd112_1 CB@23_mAd112_2 CB@23_mAd113_1 CB@23_mAd113_2 CB@23_mAd114_1 CB@23_mAd114_2 CB@23_mAd115_1 CB@23_mAd115_2 CB@23_mAd116_1 CB@23_mAd116_2 CB@23_mAd117_1 CB@23_mAd117_2 CB@23_mAd120_1 CB@23_mAd120_2 CB@23_mAd121_1 
+CB@23_mAd121_2 CB@23_mAd122_1 CB@23_mAd122_2 CB@23_mAd123_1 CB@23_mAd123_2 CB@23_mAd124_1 CB@23_mAd124_2 CB@23_mAd125_1 CB@23_mAd125_2 CB@23_mAd126_1 CB@23_mAd126_2 CB@23_mAd127_1 CB@23_mAd127_2 CB@23_mAd130_1 CB@23_mAd130_2 CB@23_mAd131_1 CB@23_mAd131_2 CB@23_mAd132_1 CB@23_mAd132_2 CB@23_mAd133_1 CB@23_mAd133_2 CB@23_mAd134_1 CB@23_mAd134_2 CB@23_mAd135_1 CB@23_mAd135_2 CB@23_mAd136_1 CB@23_mAd136_2 CB@23_mAd137_1 CB@23_mAd137_2 CB@23_mAd140_1 CB@23_mAd140_2 CB@23_mAd141_1 CB@23_mAd141_2 CB@23_mAd142_1 
+CB@23_mAd142_2 CB@23_mAd143_1 CB@23_mAd143_2 CB@23_mAd144_1 CB@23_mAd144_2 CB@23_mAd145_1 CB@23_mAd145_2 CB@23_mAd146_1 CB@23_mAd146_2 CB@23_mAd147_1 CB@23_mAd147_2 CB@23_mAd150_1 CB@23_mAd150_2 CB@23_mAd151_1 CB@23_mAd151_2 CB@23_mAd152_1 CB@23_mAd152_2 CB@23_mAd153_1 CB@23_mAd153_2 CB@23_mAd154_1 CB@23_mAd154_2 CB@23_mAd155_1 CB@23_mAd155_2 CB@23_mAd156_1 CB@23_mAd156_2 CB@23_mAd157_1 CB@23_mAd157_2 CB@23_mAd160_1 CB@23_mAd160_2 CB@23_mAd161_1 CB@23_mAd161_2 CB@23_mAd162_1 CB@23_mAd162_2 CB@23_mAd163_1 
+CB@23_mAd163_2 CB@23_mAd164_1 CB@23_mAd164_2 CB@23_mAd165_1 CB@23_mAd165_2 CB@23_mAd166_1 CB@23_mAd166_2 CB@23_mAd167_1 CB@23_mAd167_2 CB@23_mAd170_1 CB@23_mAd170_2 CB@23_mAd171_1 CB@23_mAd171_2 CB@23_mAd172_1 CB@23_mAd172_2 CB@23_mAd173_1 CB@23_mAd173_2 CB@23_mAd175_1 CB@23_mAd175_2 CB@23_mAd176_1 CB@23_mAd176_2 CB@23_mAd177_1 CB@23_mAd177_2 CB@23_mAd200_1 CB@23_mAd200_2 CB@23_mAd201_1 CB@23_mAd201_2 CB@23_mAd202_1 CB@23_mAd202_2 CB@23_mAd204_1 CB@23_mAd204_2 CB@23_mAd205_1 CB@23_mAd205_2 CB@23_mAd206_1 
+CB@23_mAd206_2 CB@23_mAd207_1 CB@23_mAd207_2 CB@23_mAd210_1 CB@23_mAd210_2 CB@23_mAd211_1 CB@23_mAd211_2 CB@23_mAd212_1 CB@23_mAd212_2 CB@23_mAd213_1 CB@23_mAd213_2 CB@23_mAd214_1 CB@23_mAd214_2 CB@23_mAd215_1 CB@23_mAd215_2 CB@23_mAd216_1 CB@23_mAd216_2 CB@23_mAd217_1 CB@23_mAd217_2 CB@23_mAd220_1 CB@23_mAd220_2 CB@23_mAd221_1 CB@23_mAd221_2 CB@23_mAd222_1 CB@23_mAd222_2 CB@23_mAd223_1 CB@23_mAd223_2 CB@23_mAd224_1 CB@23_mAd224_2 CB@23_mAd225_1 CB@23_mAd225_2 CB@23_mAd226_1 CB@23_mAd226_2 CB@23_mAd227_1 
+CB@23_mAd227_2 CB@23_mAd230_1 CB@23_mAd230_2 CB@23_mAd231_1 CB@23_mAd231_2 CB@23_mAd232_1 CB@23_mAd232_2 CB@23_mAd233_1 CB@23_mAd233_2 CB@23_mAd234_1 CB@23_mAd234_2 CB@23_mAd235_1 CB@23_mAd235_2 CB@23_mAd236_1 CB@23_mAd236_2 CB@23_mAd237_1 CB@23_mAd237_2 CB@23_mAd240_1 CB@23_mAd240_2 CB@23_mAd241_1 CB@23_mAd241_2 CB@23_mAd242_1 CB@23_mAd242_2 CB@23_mAd243_1 CB@23_mAd243_2 CB@23_mAd244_1 CB@23_mAd244_2 CB@23_mAd245_1 CB@23_mAd245_2 CB@23_mAd246_1 CB@23_mAd246_2 CB@23_mAd247_1 CB@23_mAd247_2 CB@23_mAd250_1 
+CB@23_mAd250_2 CB@23_mAd251_1 CB@23_mAd251_2 CB@23_mAd252_1 CB@23_mAd252_2 CB@23_mAd253_1 CB@23_mAd253_2 CB@23_mAd254_1 CB@23_mAd254_2 CB@23_mAd255_1 CB@23_mAd255_2 CB@23_mAd256_1 CB@23_mAd256_2 CB@23_mAd257_1 CB@23_mAd257_2 CB@23_mAd260_1 CB@23_mAd260_2 CB@23_mAd261_1 CB@23_mAd261_2 CB@23_mAd262_1 CB@23_mAd262_2 CB@23_mAd263_1 CB@23_mAd263_2 CB@23_mAd264_1 CB@23_mAd264_2 CB@23_mAd265_1 CB@23_mAd265_2 CB@23_mAd266_1 CB@23_mAd266_2 CB@23_mAd267_1 CB@23_mAd267_2 CB@23_mAd275_1 CB@23_mAd275_2 CB@23_mAd276_1 
+CB@23_mAd276_2 CB@23_mAd277_1 CB@23_mAd277_2 CB@23_mAd300_1 CB@23_mAd300_2 CB@23_mAd310_1 CB@23_mAd310_2 CB@23_mAd311_1 CB@23_mAd311_2 CB@23_mAd317_1 CB@23_mAd317_2 CB@23_mAd320_1 CB@23_mAd320_2 CB@23_mAd321_1 CB@23_mAd321_2 CB@23_mAd322_1 CB@23_mAd322_2 CB@23_mAd323_1 CB@23_mAd323_2 CB@23_mAd324_1 CB@23_mAd324_2 CB@23_mAd325_1 CB@23_mAd325_2 CB@23_mAd326_1 CB@23_mAd326_2 CB@23_mAd327_1 CB@23_mAd327_2 CB@23_mAd330_1 CB@23_mAd330_2 CB@23_mAd331_1 CB@23_mAd331_2 CB@23_mAd332_1 CB@23_mAd332_2 CB@23_mAd333_1 
+CB@23_mAd333_2 CB@23_mAd334_1 CB@23_mAd334_2 CB@23_mAd335_1 CB@23_mAd335_2 CB@23_mAd336_1 CB@23_mAd336_2 CB@23_mAd337_1 CB@23_mAd337_2 CB@23_mAd340_1 CB@23_mAd340_2 CB@23_mAd341_1 CB@23_mAd341_2 CB@23_mAd342_1 CB@23_mAd342_2 CB@23_mAd343_1 CB@23_mAd343_2 CB@23_mAd344_1 CB@23_mAd344_2 CB@23_mAd345_1 CB@23_mAd345_2 CB@23_mAd346_1 CB@23_mAd346_2 CB@23_mAd347_1 CB@23_mAd347_2 CB@23_mAd350_1 CB@23_mAd350_2 CB@23_mAd351_1 CB@23_mAd351_2 CB@23_mAd352_1 CB@23_mAd352_2 CB@23_mAd353_1 CB@23_mAd353_2 CB@23_mAd354_1 
+CB@23_mAd354_2 CB@23_mAd355_1 CB@23_mAd355_2 CB@23_mAd356_1 CB@23_mAd356_2 CB@23_mAd357_1 CB@23_mAd357_2 CB@23_mAd360_1 CB@23_mAd360_2 CB@23_mAd361_1 CB@23_mAd361_2 CB@23_mAd362_1 CB@23_mAd362_2 CB@23_mAd363_1 CB@23_mAd363_2 CB@23_mAd364_1 CB@23_mAd364_2 CB@23_mAd365_1 CB@23_mAd365_2 CB@23_mAd366_1 CB@23_mAd366_2 CB@23_mAd367_1 CB@23_mAd367_2 CB@23_mAd371_1 CB@23_mAd371_2 CB@23_mAd372_1 CB@23_mAd372_2 CB@23_mAd373_1 CB@23_mAd373_2 CB@23_mAd374_1 CB@23_mAd374_2 CB@23_mAd375_1 CB@23_mAd375_2 CB@23_mAd376_1 
+CB@23_mAd376_2 CB@23_mAd377_1 CB@23_mAd377_2 CB@23_mAd400_1 CB@23_mAd400_2 CB@23_mAd401_1 CB@23_mAd401_2 CB@23_mAd402_1 CB@23_mAd402_2 CB@23_mAd403_1 CB@23_mAd403_2 CB@23_mAd404_1 CB@23_mAd404_2 CB@23_mAd405_1 CB@23_mAd405_2 CB@23_mAd406_1 CB@23_mAd406_2 CB@23_mAd407_1 CB@23_mAd407_2 CB@23_mAd410_1 CB@23_mAd410_2 CB@23_mAd411_1 CB@23_mAd411_2 CB@23_mAd412_1 CB@23_mAd412_2 CB@23_mAd413_1 CB@23_mAd413_2 CB@23_mAd414_1 CB@23_mAd414_2 CB@23_mAd415_1 CB@23_mAd415_2 CB@23_mAd416_1 CB@23_mAd416_2 CB@23_mAd417_1 
+CB@23_mAd417_2 CB@23_mAd420_1 CB@23_mAd420_2 CB@23_mAd421_1 CB@23_mAd421_2 CB@23_mAd422_1 CB@23_mAd422_2 CB@23_mAd423_1 CB@23_mAd423_2 CB@23_mAd424_1 CB@23_mAd424_2 CB@23_mAd425_1 CB@23_mAd425_2 CB@23_mAd426_1 CB@23_mAd426_2 CB@23_mAd427_1 CB@23_mAd427_2 CB@23_mAd430_1 CB@23_mAd430_2 CB@23_mAd431_1 CB@23_mAd431_2 CB@23_mAd432_1 CB@23_mAd432_2 CB@23_mAd433_1 CB@23_mAd433_2 CB@23_mAd434_1 CB@23_mAd434_2 CB@23_mAd435_1 CB@23_mAd435_2 CB@23_mAd436_1 CB@23_mAd436_2 CB@23_mAd437_1 CB@23_mAd437_2 CB@23_mAd440_1 
+CB@23_mAd440_2 CB@23_mAd441_1 CB@23_mAd441_2 CB@23_mAd442_1 CB@23_mAd442_2 CB@23_mAd443_1 CB@23_mAd443_2 CB@23_mAd444_1 CB@23_mAd444_2 CB@23_mAd445_1 CB@23_mAd445_2 CB@23_mAd446_1 CB@23_mAd446_2 CB@23_mAd447_1 CB@23_mAd447_2 CB@23_mAd450_1 CB@23_mAd450_2 CB@23_mAd451_1 CB@23_mAd451_2 CB@23_mAd452_1 CB@23_mAd452_2 CB@23_mAd453_1 CB@23_mAd453_2 CB@23_mAd454_1 CB@23_mAd454_2 CB@23_mAd455_1 CB@23_mAd455_2 CB@23_mAd456_1 CB@23_mAd456_2 CB@23_mAd457_1 CB@23_mAd457_2 CB@23_mAd460_1 CB@23_mAd460_2 CB@23_mAd466_1 
+CB@23_mAd466_2 CB@23_mAd467_1 CB@23_mAd467_2 CB@23_mAd500_1 CB@23_mAd500_2 CB@23_mAd501_1 CB@23_mAd501_2 CB@23_mAd502_1 CB@23_mAd502_2 CB@23_mAd508_1 CB@23_mAd508_2 CB@23_mAd509_1 CB@23_mAd509_2 CB@23_mAd512_1 CB@23_mAd512_2 CB@23_mAd513_1 CB@23_mAd513_2 CB@23_mAd514_1 CB@23_mAd514_2 CB@23_mAd515_1 CB@23_mAd515_2 CB@23_mAd516_1 CB@23_mAd516_2 CB@23_mAd517_1 CB@23_mAd517_2 CB@23_mAd520_1 CB@23_mAd520_2 CB@23_mAd521_1 CB@23_mAd521_2 CB@23_mAd522_1 CB@23_mAd522_2 CB@23_mAd523_1 CB@23_mAd523_2 CB@23_mAd524_1 
+CB@23_mAd524_2 CB@23_mAd525_1 CB@23_mAd525_2 CB@23_mAd526_1 CB@23_mAd526_2 CB@23_mAd527_1 CB@23_mAd527_2 CB@23_mAd530_1 CB@23_mAd530_2 CB@23_mAd531_1 CB@23_mAd531_2 CB@23_mAd532_1 CB@23_mAd532_2 CB@23_mAd533_1 CB@23_mAd533_2 CB@23_mAd534_1 CB@23_mAd534_2 CB@23_mAd535_1 CB@23_mAd535_2 CB@23_mAd536_1 CB@23_mAd536_2 CB@23_mAd537_1 CB@23_mAd537_2 CB@23_mAd540_1 CB@23_mAd540_2 CB@23_mAd541_1 CB@23_mAd541_2 CB@23_mAd542_1 CB@23_mAd542_2 CB@23_mAd543_1 CB@23_mAd543_2 CB@23_mAd544_1 CB@23_mAd544_2 CB@23_mAd545_1 
+CB@23_mAd545_2 CB@23_mAd546_1 CB@23_mAd546_2 CB@23_mAd547_1 CB@23_mAd547_2 CB@23_mAd550_1 CB@23_mAd550_2 CB@23_mAd551_1 CB@23_mAd551_2 CB@23_mAd552_1 CB@23_mAd552_2 CB@23_mAd553_1 CB@23_mAd553_2 CB@23_mAd554_1 CB@23_mAd554_2 CB@23_mAd555_1 CB@23_mAd555_2 CB@23_mAd556_1 CB@23_mAd556_2 CB@23_mAd557_1 CB@23_mAd557_2 CB@23_mAd560_1 CB@23_mAd560_2 CB@23_mAd561_1 CB@23_mAd561_2 CB@23_mAd562_1 CB@23_mAd562_2 CB@23_mAd563_1 CB@23_mAd563_2 CB@23_mAd564_1 CB@23_mAd564_2 CB@23_mAd565_1 CB@23_mAd565_2 CB@23_mAd566_1 
+CB@23_mAd566_2 CB@23_mAd567_1 CB@23_mAd567_2 CB@23_mAd570_1 CB@23_mAd570_2 CB@23_mAd571_1 CB@23_mAd571_2 CB@23_mAd572_1 CB@23_mAd572_2 CB@23_mAd573_1 CB@23_mAd573_2 CB@23_mAd575_1 CB@23_mAd575_2 CB@23_mAd576_1 CB@23_mAd576_2 CB@23_mAd577_1 CB@23_mAd577_2 CB@23_mAd600_1 CB@23_mAd600_2 CB@23_mAd601_1 CB@23_mAd601_2 CB@23_mAd602_1 CB@23_mAd602_2 CB@23_mAd604_1 CB@23_mAd604_2 CB@23_mAd605_1 CB@23_mAd605_2 CB@23_mAd606_1 CB@23_mAd606_2 CB@23_mAd607_1 CB@23_mAd607_2 CB@23_mAd610_1 CB@23_mAd610_2 CB@23_mAd611_1 
+CB@23_mAd611_2 CB@23_mAd612_1 CB@23_mAd612_2 CB@23_mAd613_1 CB@23_mAd613_2 CB@23_mAd614_1 CB@23_mAd614_2 CB@23_mAd615_1 CB@23_mAd615_2 CB@23_mAd616_1 CB@23_mAd616_2 CB@23_mAd617_1 CB@23_mAd617_2 CB@23_mAd620_1 CB@23_mAd620_2 CB@23_mAd621_1 CB@23_mAd621_2 CB@23_mAd622_1 CB@23_mAd622_2 CB@23_mAd623_1 CB@23_mAd623_2 CB@23_mAd624_1 CB@23_mAd624_2 CB@23_mAd625_1 CB@23_mAd625_2 CB@23_mAd626_1 CB@23_mAd626_2 CB@23_mAd627_1 CB@23_mAd627_2 CB@23_mAd630_1 CB@23_mAd630_2 CB@23_mAd631_1 CB@23_mAd631_2 CB@23_mAd632_1 
+CB@23_mAd632_2 CB@23_mAd633_1 CB@23_mAd633_2 CB@23_mAd634_1 CB@23_mAd634_2 CB@23_mAd635_1 CB@23_mAd635_2 CB@23_mAd636_1 CB@23_mAd636_2 CB@23_mAd637_1 CB@23_mAd637_2 CB@23_mAd640_1 CB@23_mAd640_2 CB@23_mAd641_1 CB@23_mAd641_2 CB@23_mAd642_1 CB@23_mAd642_2 CB@23_mAd643_1 CB@23_mAd643_2 CB@23_mAd644_1 CB@23_mAd644_2 CB@23_mAd645_1 CB@23_mAd645_2 CB@23_mAd646_1 CB@23_mAd646_2 CB@23_mAd647_1 CB@23_mAd647_2 CB@23_mAd650_1 CB@23_mAd650_2 CB@23_mAd651_1 CB@23_mAd651_2 CB@23_mAd652_1 CB@23_mAd652_2 CB@23_mAd653_1 
+CB@23_mAd653_2 CB@23_mAd654_1 CB@23_mAd654_2 CB@23_mAd655_1 CB@23_mAd655_2 CB@23_mAd656_1 CB@23_mAd656_2 CB@23_mAd657_1 CB@23_mAd657_2 CB@23_mAd660_1 CB@23_mAd660_2 CB@23_mAd661_1 CB@23_mAd661_2 CB@23_mAd662_1 CB@23_mAd662_2 CB@23_mAd663_1 CB@23_mAd663_2 CB@23_mAd664_1 CB@23_mAd664_2 CB@23_mAd665_1 CB@23_mAd665_2 CB@23_mAd666_1 CB@23_mAd666_2 CB@23_mAd667_1 CB@23_mAd667_2 CB@23_mAd675_1 CB@23_mAd675_2 CB@23_mAd676_1 CB@23_mAd676_2 CB@23_mAd677_1 CB@23_mAd677_2 CB@23_mAd700_1 CB@23_mAd700_2 CB@23_mAd710_1 
+CB@23_mAd710_2 CB@23_mAd711_1 CB@23_mAd711_2 CB@23_mAd717_1 CB@23_mAd717_2 CB@23_mAd720_1 CB@23_mAd720_2 CB@23_mAd721_1 CB@23_mAd721_2 CB@23_mAd722_1 CB@23_mAd722_2 CB@23_mAd723_1 CB@23_mAd723_2 CB@23_mAd724_1 CB@23_mAd724_2 CB@23_mAd725_1 CB@23_mAd725_2 CB@23_mAd726_1 CB@23_mAd726_2 CB@23_mAd727_1 CB@23_mAd727_2 CB@23_mAd730_1 CB@23_mAd730_2 CB@23_mAd731_1 CB@23_mAd731_2 CB@23_mAd732_1 CB@23_mAd732_2 CB@23_mAd733_1 CB@23_mAd733_2 CB@23_mAd734_1 CB@23_mAd734_2 CB@23_mAd735_1 CB@23_mAd735_2 CB@23_mAd736_1 
+CB@23_mAd736_2 CB@23_mAd737_1 CB@23_mAd737_2 CB@23_mAd740_1 CB@23_mAd740_2 CB@23_mAd741_1 CB@23_mAd741_2 CB@23_mAd742_1 CB@23_mAd742_2 CB@23_mAd743_1 CB@23_mAd743_2 CB@23_mAd744_1 CB@23_mAd744_2 CB@23_mAd745_1 CB@23_mAd745_2 CB@23_mAd746_1 CB@23_mAd746_2 CB@23_mAd747_1 CB@23_mAd747_2 CB@23_mAd750_1 CB@23_mAd750_2 CB@23_mAd751_1 CB@23_mAd751_2 CB@23_mAd752_1 CB@23_mAd752_2 CB@23_mAd753_1 CB@23_mAd753_2 CB@23_mAd754_1 CB@23_mAd754_2 CB@23_mAd755_1 CB@23_mAd755_2 CB@23_mAd756_1 CB@23_mAd756_2 CB@23_mAd757_1 
+CB@23_mAd757_2 CB@23_mAd760_1 CB@23_mAd760_2 CB@23_mAd761_1 CB@23_mAd761_2 CB@23_mAd762_1 CB@23_mAd762_2 CB@23_mAd763_1 CB@23_mAd763_2 CB@23_mAd764_1 CB@23_mAd764_2 CB@23_mAd765_1 CB@23_mAd765_2 CB@23_mAd766_1 CB@23_mAd766_2 CB@23_mAd767_1 CB@23_mAd767_2 CB@23_mAd771_1 CB@23_mAd771_2 CB@23_mAd772_1 CB@23_mAd772_2 CB@23_mAd773_1 CB@23_mAd773_2 CB@23_mAd774_1 CB@23_mAd774_2 CB@23_mAd775_1 CB@23_mAd775_2 CB@23_mAd776_1 CB@23_mAd776_2 CB@23_mAd777_1 CB@23_mAd777_2 CB@23_X0 CB@23_X1 CB@23_X10 CB@23_X11 
+CB@23_X12 CB@23_X13 CB@23_X2 CB@23_X3 CB@23_X4 CB@23_X5 CB@23_X6 CB@23_X7 CB@23_X8 CB@23_X9 CB@23_Y1 CB@23_Y10 CB@23_Y11 CB@23_Y12 CB@23_Y2 CB@23_Y3 CB@23_Y4 CB@23_Y5 CB@23_Y6 CB@23_Y7 CB@23_Y8 CB@23_Y9 CB@23_Z1 CB@23_Z10 CB@23_Z11 CB@23_Z12 CB@23_Z2 CB@23_Z3 CB@23_Z4 CB@23_Z5 CB@23_Z6 CB@23_Z7 CB@23_Z8 CB@23_Z9 _5400TP094__CB
XCB@24 CB@24_K0 CB@24_K1 CB@24_K10 CB@24_K11 CB@24_K12 CB@24_K13 CB@24_K2 CB@24_K3 CB@24_K4 CB@24_K5 CB@24_K6 CB@24_K7 CB@24_K8 CB@24_K9 CB@24_mAd000_1 CB@24_mAd000_2 CB@24_mAd001_1 CB@24_mAd001_2 CB@24_mAd002_1 CB@24_mAd002_2 CB@24_mAd003_1 CB@24_mAd003_2 CB@24_mAd004_1 CB@24_mAd004_2 CB@24_mAd005_1 CB@24_mAd005_2 CB@24_mAd006_1 CB@24_mAd006_2 CB@24_mAd007_1 CB@24_mAd007_2 CB@24_mAd010_1 CB@24_mAd010_2 CB@24_mAd011_1 CB@24_mAd011_2 CB@24_mAd012_1 CB@24_mAd012_2 CB@24_mAd013_1 CB@24_mAd013_2 CB@24_mAd014_1 
+CB@24_mAd014_2 CB@24_mAd015_1 CB@24_mAd015_2 CB@24_mAd016_1 CB@24_mAd016_2 CB@24_mAd017_1 CB@24_mAd017_2 CB@24_mAd020_1 CB@24_mAd020_2 CB@24_mAd021_1 CB@24_mAd021_2 CB@24_mAd022_1 CB@24_mAd022_2 CB@24_mAd023_1 CB@24_mAd023_2 CB@24_mAd024_1 CB@24_mAd024_2 CB@24_mAd025_1 CB@24_mAd025_2 CB@24_mAd026_1 CB@24_mAd026_2 CB@24_mAd027_1 CB@24_mAd027_2 CB@24_mAd030_1 CB@24_mAd030_2 CB@24_mAd031_1 CB@24_mAd031_2 CB@24_mAd032_1 CB@24_mAd032_2 CB@24_mAd033_1 CB@24_mAd033_2 CB@24_mAd034_1 CB@24_mAd034_2 CB@24_mAd035_1 
+CB@24_mAd035_2 CB@24_mAd036_1 CB@24_mAd036_2 CB@24_mAd037_1 CB@24_mAd037_2 CB@24_mAd040_1 CB@24_mAd040_2 CB@24_mAd041_1 CB@24_mAd041_2 CB@24_mAd042_1 CB@24_mAd042_2 CB@24_mAd043_1 CB@24_mAd043_2 CB@24_mAd044_1 CB@24_mAd044_2 CB@24_mAd045_1 CB@24_mAd045_2 CB@24_mAd046_1 CB@24_mAd046_2 CB@24_mAd047_1 CB@24_mAd047_2 CB@24_mAd050_1 CB@24_mAd050_2 CB@24_mAd051_1 CB@24_mAd051_2 CB@24_mAd052_1 CB@24_mAd052_2 CB@24_mAd053_1 CB@24_mAd053_2 CB@24_mAd054_1 CB@24_mAd054_2 CB@24_mAd055_1 CB@24_mAd055_2 CB@24_mAd056_1 
+CB@24_mAd056_2 CB@24_mAd057_1 CB@24_mAd057_2 CB@24_mAd060_1 CB@24_mAd060_2 CB@24_mAd066_1 CB@24_mAd066_2 CB@24_mAd067_1 CB@24_mAd067_2 CB@24_mAd100_1 CB@24_mAd100_2 CB@24_mAd101_1 CB@24_mAd101_2 CB@24_mAd102_1 CB@24_mAd102_2 CB@24_mAd110_1 CB@24_mAd110_2 CB@24_mAd111_1 CB@24_mAd111_2 CB@24_mAd112_1 CB@24_mAd112_2 CB@24_mAd113_1 CB@24_mAd113_2 CB@24_mAd114_1 CB@24_mAd114_2 CB@24_mAd115_1 CB@24_mAd115_2 CB@24_mAd116_1 CB@24_mAd116_2 CB@24_mAd117_1 CB@24_mAd117_2 CB@24_mAd120_1 CB@24_mAd120_2 CB@24_mAd121_1 
+CB@24_mAd121_2 CB@24_mAd122_1 CB@24_mAd122_2 CB@24_mAd123_1 CB@24_mAd123_2 CB@24_mAd124_1 CB@24_mAd124_2 CB@24_mAd125_1 CB@24_mAd125_2 CB@24_mAd126_1 CB@24_mAd126_2 CB@24_mAd127_1 CB@24_mAd127_2 CB@24_mAd130_1 CB@24_mAd130_2 CB@24_mAd131_1 CB@24_mAd131_2 CB@24_mAd132_1 CB@24_mAd132_2 CB@24_mAd133_1 CB@24_mAd133_2 CB@24_mAd134_1 CB@24_mAd134_2 CB@24_mAd135_1 CB@24_mAd135_2 CB@24_mAd136_1 CB@24_mAd136_2 CB@24_mAd137_1 CB@24_mAd137_2 CB@24_mAd140_1 CB@24_mAd140_2 CB@24_mAd141_1 CB@24_mAd141_2 CB@24_mAd142_1 
+CB@24_mAd142_2 CB@24_mAd143_1 CB@24_mAd143_2 CB@24_mAd144_1 CB@24_mAd144_2 CB@24_mAd145_1 CB@24_mAd145_2 CB@24_mAd146_1 CB@24_mAd146_2 CB@24_mAd147_1 CB@24_mAd147_2 CB@24_mAd150_1 CB@24_mAd150_2 CB@24_mAd151_1 CB@24_mAd151_2 CB@24_mAd152_1 CB@24_mAd152_2 CB@24_mAd153_1 CB@24_mAd153_2 CB@24_mAd154_1 CB@24_mAd154_2 CB@24_mAd155_1 CB@24_mAd155_2 CB@24_mAd156_1 CB@24_mAd156_2 CB@24_mAd157_1 CB@24_mAd157_2 CB@24_mAd160_1 CB@24_mAd160_2 CB@24_mAd161_1 CB@24_mAd161_2 CB@24_mAd162_1 CB@24_mAd162_2 CB@24_mAd163_1 
+CB@24_mAd163_2 CB@24_mAd164_1 CB@24_mAd164_2 CB@24_mAd165_1 CB@24_mAd165_2 CB@24_mAd166_1 CB@24_mAd166_2 CB@24_mAd167_1 CB@24_mAd167_2 CB@24_mAd170_1 CB@24_mAd170_2 CB@24_mAd171_1 CB@24_mAd171_2 CB@24_mAd172_1 CB@24_mAd172_2 CB@24_mAd173_1 CB@24_mAd173_2 CB@24_mAd175_1 CB@24_mAd175_2 CB@24_mAd176_1 CB@24_mAd176_2 CB@24_mAd177_1 CB@24_mAd177_2 CB@24_mAd200_1 CB@24_mAd200_2 CB@24_mAd201_1 CB@24_mAd201_2 CB@24_mAd202_1 CB@24_mAd202_2 CB@24_mAd204_1 CB@24_mAd204_2 CB@24_mAd205_1 CB@24_mAd205_2 CB@24_mAd206_1 
+CB@24_mAd206_2 CB@24_mAd207_1 CB@24_mAd207_2 CB@24_mAd210_1 CB@24_mAd210_2 CB@24_mAd211_1 CB@24_mAd211_2 CB@24_mAd212_1 CB@24_mAd212_2 CB@24_mAd213_1 CB@24_mAd213_2 CB@24_mAd214_1 CB@24_mAd214_2 CB@24_mAd215_1 CB@24_mAd215_2 CB@24_mAd216_1 CB@24_mAd216_2 CB@24_mAd217_1 CB@24_mAd217_2 CB@24_mAd220_1 CB@24_mAd220_2 CB@24_mAd221_1 CB@24_mAd221_2 CB@24_mAd222_1 CB@24_mAd222_2 CB@24_mAd223_1 CB@24_mAd223_2 CB@24_mAd224_1 CB@24_mAd224_2 CB@24_mAd225_1 CB@24_mAd225_2 CB@24_mAd226_1 CB@24_mAd226_2 CB@24_mAd227_1 
+CB@24_mAd227_2 CB@24_mAd230_1 CB@24_mAd230_2 CB@24_mAd231_1 CB@24_mAd231_2 CB@24_mAd232_1 CB@24_mAd232_2 CB@24_mAd233_1 CB@24_mAd233_2 CB@24_mAd234_1 CB@24_mAd234_2 CB@24_mAd235_1 CB@24_mAd235_2 CB@24_mAd236_1 CB@24_mAd236_2 CB@24_mAd237_1 CB@24_mAd237_2 CB@24_mAd240_1 CB@24_mAd240_2 CB@24_mAd241_1 CB@24_mAd241_2 CB@24_mAd242_1 CB@24_mAd242_2 CB@24_mAd243_1 CB@24_mAd243_2 CB@24_mAd244_1 CB@24_mAd244_2 CB@24_mAd245_1 CB@24_mAd245_2 CB@24_mAd246_1 CB@24_mAd246_2 CB@24_mAd247_1 CB@24_mAd247_2 CB@24_mAd250_1 
+CB@24_mAd250_2 CB@24_mAd251_1 CB@24_mAd251_2 CB@24_mAd252_1 CB@24_mAd252_2 CB@24_mAd253_1 CB@24_mAd253_2 CB@24_mAd254_1 CB@24_mAd254_2 CB@24_mAd255_1 CB@24_mAd255_2 CB@24_mAd256_1 CB@24_mAd256_2 CB@24_mAd257_1 CB@24_mAd257_2 CB@24_mAd260_1 CB@24_mAd260_2 CB@24_mAd261_1 CB@24_mAd261_2 CB@24_mAd262_1 CB@24_mAd262_2 CB@24_mAd263_1 CB@24_mAd263_2 CB@24_mAd264_1 CB@24_mAd264_2 CB@24_mAd265_1 CB@24_mAd265_2 CB@24_mAd266_1 CB@24_mAd266_2 CB@24_mAd267_1 CB@24_mAd267_2 CB@24_mAd275_1 CB@24_mAd275_2 CB@24_mAd276_1 
+CB@24_mAd276_2 CB@24_mAd277_1 CB@24_mAd277_2 CB@24_mAd300_1 CB@24_mAd300_2 CB@24_mAd310_1 CB@24_mAd310_2 CB@24_mAd311_1 CB@24_mAd311_2 CB@24_mAd317_1 CB@24_mAd317_2 CB@24_mAd320_1 CB@24_mAd320_2 CB@24_mAd321_1 CB@24_mAd321_2 CB@24_mAd322_1 CB@24_mAd322_2 CB@24_mAd323_1 CB@24_mAd323_2 CB@24_mAd324_1 CB@24_mAd324_2 CB@24_mAd325_1 CB@24_mAd325_2 CB@24_mAd326_1 CB@24_mAd326_2 CB@24_mAd327_1 CB@24_mAd327_2 CB@24_mAd330_1 CB@24_mAd330_2 CB@24_mAd331_1 CB@24_mAd331_2 CB@24_mAd332_1 CB@24_mAd332_2 CB@24_mAd333_1 
+CB@24_mAd333_2 CB@24_mAd334_1 CB@24_mAd334_2 CB@24_mAd335_1 CB@24_mAd335_2 CB@24_mAd336_1 CB@24_mAd336_2 CB@24_mAd337_1 CB@24_mAd337_2 CB@24_mAd340_1 CB@24_mAd340_2 CB@24_mAd341_1 CB@24_mAd341_2 CB@24_mAd342_1 CB@24_mAd342_2 CB@24_mAd343_1 CB@24_mAd343_2 CB@24_mAd344_1 CB@24_mAd344_2 CB@24_mAd345_1 CB@24_mAd345_2 CB@24_mAd346_1 CB@24_mAd346_2 CB@24_mAd347_1 CB@24_mAd347_2 CB@24_mAd350_1 CB@24_mAd350_2 CB@24_mAd351_1 CB@24_mAd351_2 CB@24_mAd352_1 CB@24_mAd352_2 CB@24_mAd353_1 CB@24_mAd353_2 CB@24_mAd354_1 
+CB@24_mAd354_2 CB@24_mAd355_1 CB@24_mAd355_2 CB@24_mAd356_1 CB@24_mAd356_2 CB@24_mAd357_1 CB@24_mAd357_2 CB@24_mAd360_1 CB@24_mAd360_2 CB@24_mAd361_1 CB@24_mAd361_2 CB@24_mAd362_1 CB@24_mAd362_2 CB@24_mAd363_1 CB@24_mAd363_2 CB@24_mAd364_1 CB@24_mAd364_2 CB@24_mAd365_1 CB@24_mAd365_2 CB@24_mAd366_1 CB@24_mAd366_2 CB@24_mAd367_1 CB@24_mAd367_2 CB@24_mAd371_1 CB@24_mAd371_2 CB@24_mAd372_1 CB@24_mAd372_2 CB@24_mAd373_1 CB@24_mAd373_2 CB@24_mAd374_1 CB@24_mAd374_2 CB@24_mAd375_1 CB@24_mAd375_2 CB@24_mAd376_1 
+CB@24_mAd376_2 CB@24_mAd377_1 CB@24_mAd377_2 CB@24_mAd400_1 CB@24_mAd400_2 CB@24_mAd401_1 CB@24_mAd401_2 CB@24_mAd402_1 CB@24_mAd402_2 CB@24_mAd403_1 CB@24_mAd403_2 CB@24_mAd404_1 CB@24_mAd404_2 CB@24_mAd405_1 CB@24_mAd405_2 CB@24_mAd406_1 CB@24_mAd406_2 CB@24_mAd407_1 CB@24_mAd407_2 CB@24_mAd410_1 CB@24_mAd410_2 CB@24_mAd411_1 CB@24_mAd411_2 CB@24_mAd412_1 CB@24_mAd412_2 CB@24_mAd413_1 CB@24_mAd413_2 CB@24_mAd414_1 CB@24_mAd414_2 CB@24_mAd415_1 CB@24_mAd415_2 CB@24_mAd416_1 CB@24_mAd416_2 CB@24_mAd417_1 
+CB@24_mAd417_2 CB@24_mAd420_1 CB@24_mAd420_2 CB@24_mAd421_1 CB@24_mAd421_2 CB@24_mAd422_1 CB@24_mAd422_2 CB@24_mAd423_1 CB@24_mAd423_2 CB@24_mAd424_1 CB@24_mAd424_2 CB@24_mAd425_1 CB@24_mAd425_2 CB@24_mAd426_1 CB@24_mAd426_2 CB@24_mAd427_1 CB@24_mAd427_2 CB@24_mAd430_1 CB@24_mAd430_2 CB@24_mAd431_1 CB@24_mAd431_2 CB@24_mAd432_1 CB@24_mAd432_2 CB@24_mAd433_1 CB@24_mAd433_2 CB@24_mAd434_1 CB@24_mAd434_2 CB@24_mAd435_1 CB@24_mAd435_2 CB@24_mAd436_1 CB@24_mAd436_2 CB@24_mAd437_1 CB@24_mAd437_2 CB@24_mAd440_1 
+CB@24_mAd440_2 CB@24_mAd441_1 CB@24_mAd441_2 CB@24_mAd442_1 CB@24_mAd442_2 CB@24_mAd443_1 CB@24_mAd443_2 CB@24_mAd444_1 CB@24_mAd444_2 CB@24_mAd445_1 CB@24_mAd445_2 CB@24_mAd446_1 CB@24_mAd446_2 CB@24_mAd447_1 CB@24_mAd447_2 CB@24_mAd450_1 CB@24_mAd450_2 CB@24_mAd451_1 CB@24_mAd451_2 CB@24_mAd452_1 CB@24_mAd452_2 CB@24_mAd453_1 CB@24_mAd453_2 CB@24_mAd454_1 CB@24_mAd454_2 CB@24_mAd455_1 CB@24_mAd455_2 CB@24_mAd456_1 CB@24_mAd456_2 CB@24_mAd457_1 CB@24_mAd457_2 CB@24_mAd460_1 CB@24_mAd460_2 CB@24_mAd466_1 
+CB@24_mAd466_2 CB@24_mAd467_1 CB@24_mAd467_2 CB@24_mAd500_1 CB@24_mAd500_2 CB@24_mAd501_1 CB@24_mAd501_2 CB@24_mAd502_1 CB@24_mAd502_2 CB@24_mAd508_1 CB@24_mAd508_2 CB@24_mAd509_1 CB@24_mAd509_2 CB@24_mAd512_1 CB@24_mAd512_2 CB@24_mAd513_1 CB@24_mAd513_2 CB@24_mAd514_1 CB@24_mAd514_2 CB@24_mAd515_1 CB@24_mAd515_2 CB@24_mAd516_1 CB@24_mAd516_2 CB@24_mAd517_1 CB@24_mAd517_2 CB@24_mAd520_1 CB@24_mAd520_2 CB@24_mAd521_1 CB@24_mAd521_2 CB@24_mAd522_1 CB@24_mAd522_2 CB@24_mAd523_1 CB@24_mAd523_2 CB@24_mAd524_1 
+CB@24_mAd524_2 CB@24_mAd525_1 CB@24_mAd525_2 CB@24_mAd526_1 CB@24_mAd526_2 CB@24_mAd527_1 CB@24_mAd527_2 CB@24_mAd530_1 CB@24_mAd530_2 CB@24_mAd531_1 CB@24_mAd531_2 CB@24_mAd532_1 CB@24_mAd532_2 CB@24_mAd533_1 CB@24_mAd533_2 CB@24_mAd534_1 CB@24_mAd534_2 CB@24_mAd535_1 CB@24_mAd535_2 CB@24_mAd536_1 CB@24_mAd536_2 CB@24_mAd537_1 CB@24_mAd537_2 CB@24_mAd540_1 CB@24_mAd540_2 CB@24_mAd541_1 CB@24_mAd541_2 CB@24_mAd542_1 CB@24_mAd542_2 CB@24_mAd543_1 CB@24_mAd543_2 CB@24_mAd544_1 CB@24_mAd544_2 CB@24_mAd545_1 
+CB@24_mAd545_2 CB@24_mAd546_1 CB@24_mAd546_2 CB@24_mAd547_1 CB@24_mAd547_2 CB@24_mAd550_1 CB@24_mAd550_2 CB@24_mAd551_1 CB@24_mAd551_2 CB@24_mAd552_1 CB@24_mAd552_2 CB@24_mAd553_1 CB@24_mAd553_2 CB@24_mAd554_1 CB@24_mAd554_2 CB@24_mAd555_1 CB@24_mAd555_2 CB@24_mAd556_1 CB@24_mAd556_2 CB@24_mAd557_1 CB@24_mAd557_2 CB@24_mAd560_1 CB@24_mAd560_2 CB@24_mAd561_1 CB@24_mAd561_2 CB@24_mAd562_1 CB@24_mAd562_2 CB@24_mAd563_1 CB@24_mAd563_2 CB@24_mAd564_1 CB@24_mAd564_2 CB@24_mAd565_1 CB@24_mAd565_2 CB@24_mAd566_1 
+CB@24_mAd566_2 CB@24_mAd567_1 CB@24_mAd567_2 CB@24_mAd570_1 CB@24_mAd570_2 CB@24_mAd571_1 CB@24_mAd571_2 CB@24_mAd572_1 CB@24_mAd572_2 CB@24_mAd573_1 CB@24_mAd573_2 CB@24_mAd575_1 CB@24_mAd575_2 CB@24_mAd576_1 CB@24_mAd576_2 CB@24_mAd577_1 CB@24_mAd577_2 CB@24_mAd600_1 CB@24_mAd600_2 CB@24_mAd601_1 CB@24_mAd601_2 CB@24_mAd602_1 CB@24_mAd602_2 CB@24_mAd604_1 CB@24_mAd604_2 CB@24_mAd605_1 CB@24_mAd605_2 CB@24_mAd606_1 CB@24_mAd606_2 CB@24_mAd607_1 CB@24_mAd607_2 CB@24_mAd610_1 CB@24_mAd610_2 CB@24_mAd611_1 
+CB@24_mAd611_2 CB@24_mAd612_1 CB@24_mAd612_2 CB@24_mAd613_1 CB@24_mAd613_2 CB@24_mAd614_1 CB@24_mAd614_2 CB@24_mAd615_1 CB@24_mAd615_2 CB@24_mAd616_1 CB@24_mAd616_2 CB@24_mAd617_1 CB@24_mAd617_2 CB@24_mAd620_1 CB@24_mAd620_2 CB@24_mAd621_1 CB@24_mAd621_2 CB@24_mAd622_1 CB@24_mAd622_2 CB@24_mAd623_1 CB@24_mAd623_2 CB@24_mAd624_1 CB@24_mAd624_2 CB@24_mAd625_1 CB@24_mAd625_2 CB@24_mAd626_1 CB@24_mAd626_2 CB@24_mAd627_1 CB@24_mAd627_2 CB@24_mAd630_1 CB@24_mAd630_2 CB@24_mAd631_1 CB@24_mAd631_2 CB@24_mAd632_1 
+CB@24_mAd632_2 CB@24_mAd633_1 CB@24_mAd633_2 CB@24_mAd634_1 CB@24_mAd634_2 CB@24_mAd635_1 CB@24_mAd635_2 CB@24_mAd636_1 CB@24_mAd636_2 CB@24_mAd637_1 CB@24_mAd637_2 CB@24_mAd640_1 CB@24_mAd640_2 CB@24_mAd641_1 CB@24_mAd641_2 CB@24_mAd642_1 CB@24_mAd642_2 CB@24_mAd643_1 CB@24_mAd643_2 CB@24_mAd644_1 CB@24_mAd644_2 CB@24_mAd645_1 CB@24_mAd645_2 CB@24_mAd646_1 CB@24_mAd646_2 CB@24_mAd647_1 CB@24_mAd647_2 CB@24_mAd650_1 CB@24_mAd650_2 CB@24_mAd651_1 CB@24_mAd651_2 CB@24_mAd652_1 CB@24_mAd652_2 CB@24_mAd653_1 
+CB@24_mAd653_2 CB@24_mAd654_1 CB@24_mAd654_2 CB@24_mAd655_1 CB@24_mAd655_2 CB@24_mAd656_1 CB@24_mAd656_2 CB@24_mAd657_1 CB@24_mAd657_2 CB@24_mAd660_1 CB@24_mAd660_2 CB@24_mAd661_1 CB@24_mAd661_2 CB@24_mAd662_1 CB@24_mAd662_2 CB@24_mAd663_1 CB@24_mAd663_2 CB@24_mAd664_1 CB@24_mAd664_2 CB@24_mAd665_1 CB@24_mAd665_2 CB@24_mAd666_1 CB@24_mAd666_2 CB@24_mAd667_1 CB@24_mAd667_2 CB@24_mAd675_1 CB@24_mAd675_2 CB@24_mAd676_1 CB@24_mAd676_2 CB@24_mAd677_1 CB@24_mAd677_2 CB@24_mAd700_1 CB@24_mAd700_2 CB@24_mAd710_1 
+CB@24_mAd710_2 CB@24_mAd711_1 CB@24_mAd711_2 CB@24_mAd717_1 CB@24_mAd717_2 CB@24_mAd720_1 CB@24_mAd720_2 CB@24_mAd721_1 CB@24_mAd721_2 CB@24_mAd722_1 CB@24_mAd722_2 CB@24_mAd723_1 CB@24_mAd723_2 CB@24_mAd724_1 CB@24_mAd724_2 CB@24_mAd725_1 CB@24_mAd725_2 CB@24_mAd726_1 CB@24_mAd726_2 CB@24_mAd727_1 CB@24_mAd727_2 CB@24_mAd730_1 CB@24_mAd730_2 CB@24_mAd731_1 CB@24_mAd731_2 CB@24_mAd732_1 CB@24_mAd732_2 CB@24_mAd733_1 CB@24_mAd733_2 CB@24_mAd734_1 CB@24_mAd734_2 CB@24_mAd735_1 CB@24_mAd735_2 CB@24_mAd736_1 
+CB@24_mAd736_2 CB@24_mAd737_1 CB@24_mAd737_2 CB@24_mAd740_1 CB@24_mAd740_2 CB@24_mAd741_1 CB@24_mAd741_2 CB@24_mAd742_1 CB@24_mAd742_2 CB@24_mAd743_1 CB@24_mAd743_2 CB@24_mAd744_1 CB@24_mAd744_2 CB@24_mAd745_1 CB@24_mAd745_2 CB@24_mAd746_1 CB@24_mAd746_2 CB@24_mAd747_1 CB@24_mAd747_2 CB@24_mAd750_1 CB@24_mAd750_2 CB@24_mAd751_1 CB@24_mAd751_2 CB@24_mAd752_1 CB@24_mAd752_2 CB@24_mAd753_1 CB@24_mAd753_2 CB@24_mAd754_1 CB@24_mAd754_2 CB@24_mAd755_1 CB@24_mAd755_2 CB@24_mAd756_1 CB@24_mAd756_2 CB@24_mAd757_1 
+CB@24_mAd757_2 CB@24_mAd760_1 CB@24_mAd760_2 CB@24_mAd761_1 CB@24_mAd761_2 CB@24_mAd762_1 CB@24_mAd762_2 CB@24_mAd763_1 CB@24_mAd763_2 CB@24_mAd764_1 CB@24_mAd764_2 CB@24_mAd765_1 CB@24_mAd765_2 CB@24_mAd766_1 CB@24_mAd766_2 CB@24_mAd767_1 CB@24_mAd767_2 CB@24_mAd771_1 CB@24_mAd771_2 CB@24_mAd772_1 CB@24_mAd772_2 CB@24_mAd773_1 CB@24_mAd773_2 CB@24_mAd774_1 CB@24_mAd774_2 CB@24_mAd775_1 CB@24_mAd775_2 CB@24_mAd776_1 CB@24_mAd776_2 CB@24_mAd777_1 CB@24_mAd777_2 CB@24_X0 CB@24_X1 CB@24_X10 CB@24_X11 
+CB@24_X12 CB@24_X13 CB@24_X2 CB@24_X3 CB@24_X4 CB@24_X5 CB@24_X6 CB@24_X7 CB@24_X8 CB@24_X9 CB@24_Y1 CB@24_Y10 CB@24_Y11 CB@24_Y12 CB@24_Y2 CB@24_Y3 CB@24_Y4 CB@24_Y5 CB@24_Y6 CB@24_Y7 CB@24_Y8 CB@24_Y9 CB@24_Z1 CB@24_Z10 CB@24_Z11 CB@24_Z12 CB@24_Z2 CB@24_Z3 CB@24_Z4 CB@24_Z5 CB@24_Z6 CB@24_Z7 CB@24_Z8 CB@24_Z9 _5400TP094__CB
XCB@25 CB@25_K0 CB@25_K1 CB@25_K10 CB@25_K11 CB@25_K12 CB@25_K13 CB@25_K2 CB@25_K3 CB@25_K4 CB@25_K5 CB@25_K6 CB@25_K7 CB@25_K8 CB@25_K9 CB@25_mAd000_1 CB@25_mAd000_2 CB@25_mAd001_1 CB@25_mAd001_2 CB@25_mAd002_1 CB@25_mAd002_2 CB@25_mAd003_1 CB@25_mAd003_2 CB@25_mAd004_1 CB@25_mAd004_2 CB@25_mAd005_1 CB@25_mAd005_2 CB@25_mAd006_1 CB@25_mAd006_2 CB@25_mAd007_1 CB@25_mAd007_2 CB@25_mAd010_1 CB@25_mAd010_2 CB@25_mAd011_1 CB@25_mAd011_2 CB@25_mAd012_1 CB@25_mAd012_2 CB@25_mAd013_1 CB@25_mAd013_2 CB@25_mAd014_1 
+CB@25_mAd014_2 CB@25_mAd015_1 CB@25_mAd015_2 CB@25_mAd016_1 CB@25_mAd016_2 CB@25_mAd017_1 CB@25_mAd017_2 CB@25_mAd020_1 CB@25_mAd020_2 CB@25_mAd021_1 CB@25_mAd021_2 CB@25_mAd022_1 CB@25_mAd022_2 CB@25_mAd023_1 CB@25_mAd023_2 CB@25_mAd024_1 CB@25_mAd024_2 CB@25_mAd025_1 CB@25_mAd025_2 CB@25_mAd026_1 CB@25_mAd026_2 CB@25_mAd027_1 CB@25_mAd027_2 CB@25_mAd030_1 CB@25_mAd030_2 CB@25_mAd031_1 CB@25_mAd031_2 CB@25_mAd032_1 CB@25_mAd032_2 CB@25_mAd033_1 CB@25_mAd033_2 CB@25_mAd034_1 CB@25_mAd034_2 CB@25_mAd035_1 
+CB@25_mAd035_2 CB@25_mAd036_1 CB@25_mAd036_2 CB@25_mAd037_1 CB@25_mAd037_2 CB@25_mAd040_1 CB@25_mAd040_2 CB@25_mAd041_1 CB@25_mAd041_2 CB@25_mAd042_1 CB@25_mAd042_2 CB@25_mAd043_1 CB@25_mAd043_2 CB@25_mAd044_1 CB@25_mAd044_2 CB@25_mAd045_1 CB@25_mAd045_2 CB@25_mAd046_1 CB@25_mAd046_2 CB@25_mAd047_1 CB@25_mAd047_2 CB@25_mAd050_1 CB@25_mAd050_2 CB@25_mAd051_1 CB@25_mAd051_2 CB@25_mAd052_1 CB@25_mAd052_2 CB@25_mAd053_1 CB@25_mAd053_2 CB@25_mAd054_1 CB@25_mAd054_2 CB@25_mAd055_1 CB@25_mAd055_2 CB@25_mAd056_1 
+CB@25_mAd056_2 CB@25_mAd057_1 CB@25_mAd057_2 CB@25_mAd060_1 CB@25_mAd060_2 CB@25_mAd066_1 CB@25_mAd066_2 CB@25_mAd067_1 CB@25_mAd067_2 CB@25_mAd100_1 CB@25_mAd100_2 CB@25_mAd101_1 CB@25_mAd101_2 CB@25_mAd102_1 CB@25_mAd102_2 CB@25_mAd110_1 CB@25_mAd110_2 CB@25_mAd111_1 CB@25_mAd111_2 CB@25_mAd112_1 CB@25_mAd112_2 CB@25_mAd113_1 CB@25_mAd113_2 CB@25_mAd114_1 CB@25_mAd114_2 CB@25_mAd115_1 CB@25_mAd115_2 CB@25_mAd116_1 CB@25_mAd116_2 CB@25_mAd117_1 CB@25_mAd117_2 CB@25_mAd120_1 CB@25_mAd120_2 CB@25_mAd121_1 
+CB@25_mAd121_2 CB@25_mAd122_1 CB@25_mAd122_2 CB@25_mAd123_1 CB@25_mAd123_2 CB@25_mAd124_1 CB@25_mAd124_2 CB@25_mAd125_1 CB@25_mAd125_2 CB@25_mAd126_1 CB@25_mAd126_2 CB@25_mAd127_1 CB@25_mAd127_2 CB@25_mAd130_1 CB@25_mAd130_2 CB@25_mAd131_1 CB@25_mAd131_2 CB@25_mAd132_1 CB@25_mAd132_2 CB@25_mAd133_1 CB@25_mAd133_2 CB@25_mAd134_1 CB@25_mAd134_2 CB@25_mAd135_1 CB@25_mAd135_2 CB@25_mAd136_1 CB@25_mAd136_2 CB@25_mAd137_1 CB@25_mAd137_2 CB@25_mAd140_1 CB@25_mAd140_2 CB@25_mAd141_1 CB@25_mAd141_2 CB@25_mAd142_1 
+CB@25_mAd142_2 CB@25_mAd143_1 CB@25_mAd143_2 CB@25_mAd144_1 CB@25_mAd144_2 CB@25_mAd145_1 CB@25_mAd145_2 CB@25_mAd146_1 CB@25_mAd146_2 CB@25_mAd147_1 CB@25_mAd147_2 CB@25_mAd150_1 CB@25_mAd150_2 CB@25_mAd151_1 CB@25_mAd151_2 CB@25_mAd152_1 CB@25_mAd152_2 CB@25_mAd153_1 CB@25_mAd153_2 CB@25_mAd154_1 CB@25_mAd154_2 CB@25_mAd155_1 CB@25_mAd155_2 CB@25_mAd156_1 CB@25_mAd156_2 CB@25_mAd157_1 CB@25_mAd157_2 CB@25_mAd160_1 CB@25_mAd160_2 CB@25_mAd161_1 CB@25_mAd161_2 CB@25_mAd162_1 CB@25_mAd162_2 CB@25_mAd163_1 
+CB@25_mAd163_2 CB@25_mAd164_1 CB@25_mAd164_2 CB@25_mAd165_1 CB@25_mAd165_2 CB@25_mAd166_1 CB@25_mAd166_2 CB@25_mAd167_1 CB@25_mAd167_2 CB@25_mAd170_1 CB@25_mAd170_2 CB@25_mAd171_1 CB@25_mAd171_2 CB@25_mAd172_1 CB@25_mAd172_2 CB@25_mAd173_1 CB@25_mAd173_2 CB@25_mAd175_1 CB@25_mAd175_2 CB@25_mAd176_1 CB@25_mAd176_2 CB@25_mAd177_1 CB@25_mAd177_2 CB@25_mAd200_1 CB@25_mAd200_2 CB@25_mAd201_1 CB@25_mAd201_2 CB@25_mAd202_1 CB@25_mAd202_2 CB@25_mAd204_1 CB@25_mAd204_2 CB@25_mAd205_1 CB@25_mAd205_2 CB@25_mAd206_1 
+CB@25_mAd206_2 CB@25_mAd207_1 CB@25_mAd207_2 CB@25_mAd210_1 CB@25_mAd210_2 CB@25_mAd211_1 CB@25_mAd211_2 CB@25_mAd212_1 CB@25_mAd212_2 CB@25_mAd213_1 CB@25_mAd213_2 CB@25_mAd214_1 CB@25_mAd214_2 CB@25_mAd215_1 CB@25_mAd215_2 CB@25_mAd216_1 CB@25_mAd216_2 CB@25_mAd217_1 CB@25_mAd217_2 CB@25_mAd220_1 CB@25_mAd220_2 CB@25_mAd221_1 CB@25_mAd221_2 CB@25_mAd222_1 CB@25_mAd222_2 CB@25_mAd223_1 CB@25_mAd223_2 CB@25_mAd224_1 CB@25_mAd224_2 CB@25_mAd225_1 CB@25_mAd225_2 CB@25_mAd226_1 CB@25_mAd226_2 CB@25_mAd227_1 
+CB@25_mAd227_2 CB@25_mAd230_1 CB@25_mAd230_2 CB@25_mAd231_1 CB@25_mAd231_2 CB@25_mAd232_1 CB@25_mAd232_2 CB@25_mAd233_1 CB@25_mAd233_2 CB@25_mAd234_1 CB@25_mAd234_2 CB@25_mAd235_1 CB@25_mAd235_2 CB@25_mAd236_1 CB@25_mAd236_2 CB@25_mAd237_1 CB@25_mAd237_2 CB@25_mAd240_1 CB@25_mAd240_2 CB@25_mAd241_1 CB@25_mAd241_2 CB@25_mAd242_1 CB@25_mAd242_2 CB@25_mAd243_1 CB@25_mAd243_2 CB@25_mAd244_1 CB@25_mAd244_2 CB@25_mAd245_1 CB@25_mAd245_2 CB@25_mAd246_1 CB@25_mAd246_2 CB@25_mAd247_1 CB@25_mAd247_2 CB@25_mAd250_1 
+CB@25_mAd250_2 CB@25_mAd251_1 CB@25_mAd251_2 CB@25_mAd252_1 CB@25_mAd252_2 CB@25_mAd253_1 CB@25_mAd253_2 CB@25_mAd254_1 CB@25_mAd254_2 CB@25_mAd255_1 CB@25_mAd255_2 CB@25_mAd256_1 CB@25_mAd256_2 CB@25_mAd257_1 CB@25_mAd257_2 CB@25_mAd260_1 CB@25_mAd260_2 CB@25_mAd261_1 CB@25_mAd261_2 CB@25_mAd262_1 CB@25_mAd262_2 CB@25_mAd263_1 CB@25_mAd263_2 CB@25_mAd264_1 CB@25_mAd264_2 CB@25_mAd265_1 CB@25_mAd265_2 CB@25_mAd266_1 CB@25_mAd266_2 CB@25_mAd267_1 CB@25_mAd267_2 CB@25_mAd275_1 CB@25_mAd275_2 CB@25_mAd276_1 
+CB@25_mAd276_2 CB@25_mAd277_1 CB@25_mAd277_2 CB@25_mAd300_1 CB@25_mAd300_2 CB@25_mAd310_1 CB@25_mAd310_2 CB@25_mAd311_1 CB@25_mAd311_2 CB@25_mAd317_1 CB@25_mAd317_2 CB@25_mAd320_1 CB@25_mAd320_2 CB@25_mAd321_1 CB@25_mAd321_2 CB@25_mAd322_1 CB@25_mAd322_2 CB@25_mAd323_1 CB@25_mAd323_2 CB@25_mAd324_1 CB@25_mAd324_2 CB@25_mAd325_1 CB@25_mAd325_2 CB@25_mAd326_1 CB@25_mAd326_2 CB@25_mAd327_1 CB@25_mAd327_2 CB@25_mAd330_1 CB@25_mAd330_2 CB@25_mAd331_1 CB@25_mAd331_2 CB@25_mAd332_1 CB@25_mAd332_2 CB@25_mAd333_1 
+CB@25_mAd333_2 CB@25_mAd334_1 CB@25_mAd334_2 CB@25_mAd335_1 CB@25_mAd335_2 CB@25_mAd336_1 CB@25_mAd336_2 CB@25_mAd337_1 CB@25_mAd337_2 CB@25_mAd340_1 CB@25_mAd340_2 CB@25_mAd341_1 CB@25_mAd341_2 CB@25_mAd342_1 CB@25_mAd342_2 CB@25_mAd343_1 CB@25_mAd343_2 CB@25_mAd344_1 CB@25_mAd344_2 CB@25_mAd345_1 CB@25_mAd345_2 CB@25_mAd346_1 CB@25_mAd346_2 CB@25_mAd347_1 CB@25_mAd347_2 CB@25_mAd350_1 CB@25_mAd350_2 CB@25_mAd351_1 CB@25_mAd351_2 CB@25_mAd352_1 CB@25_mAd352_2 CB@25_mAd353_1 CB@25_mAd353_2 CB@25_mAd354_1 
+CB@25_mAd354_2 CB@25_mAd355_1 CB@25_mAd355_2 CB@25_mAd356_1 CB@25_mAd356_2 CB@25_mAd357_1 CB@25_mAd357_2 CB@25_mAd360_1 CB@25_mAd360_2 CB@25_mAd361_1 CB@25_mAd361_2 CB@25_mAd362_1 CB@25_mAd362_2 CB@25_mAd363_1 CB@25_mAd363_2 CB@25_mAd364_1 CB@25_mAd364_2 CB@25_mAd365_1 CB@25_mAd365_2 CB@25_mAd366_1 CB@25_mAd366_2 CB@25_mAd367_1 CB@25_mAd367_2 CB@25_mAd371_1 CB@25_mAd371_2 CB@25_mAd372_1 CB@25_mAd372_2 CB@25_mAd373_1 CB@25_mAd373_2 CB@25_mAd374_1 CB@25_mAd374_2 CB@25_mAd375_1 CB@25_mAd375_2 CB@25_mAd376_1 
+CB@25_mAd376_2 CB@25_mAd377_1 CB@25_mAd377_2 CB@25_mAd400_1 CB@25_mAd400_2 CB@25_mAd401_1 CB@25_mAd401_2 CB@25_mAd402_1 CB@25_mAd402_2 CB@25_mAd403_1 CB@25_mAd403_2 CB@25_mAd404_1 CB@25_mAd404_2 CB@25_mAd405_1 CB@25_mAd405_2 CB@25_mAd406_1 CB@25_mAd406_2 CB@25_mAd407_1 CB@25_mAd407_2 CB@25_mAd410_1 CB@25_mAd410_2 CB@25_mAd411_1 CB@25_mAd411_2 CB@25_mAd412_1 CB@25_mAd412_2 CB@25_mAd413_1 CB@25_mAd413_2 CB@25_mAd414_1 CB@25_mAd414_2 CB@25_mAd415_1 CB@25_mAd415_2 CB@25_mAd416_1 CB@25_mAd416_2 CB@25_mAd417_1 
+CB@25_mAd417_2 CB@25_mAd420_1 CB@25_mAd420_2 CB@25_mAd421_1 CB@25_mAd421_2 CB@25_mAd422_1 CB@25_mAd422_2 CB@25_mAd423_1 CB@25_mAd423_2 CB@25_mAd424_1 CB@25_mAd424_2 CB@25_mAd425_1 CB@25_mAd425_2 CB@25_mAd426_1 CB@25_mAd426_2 CB@25_mAd427_1 CB@25_mAd427_2 CB@25_mAd430_1 CB@25_mAd430_2 CB@25_mAd431_1 CB@25_mAd431_2 CB@25_mAd432_1 CB@25_mAd432_2 CB@25_mAd433_1 CB@25_mAd433_2 CB@25_mAd434_1 CB@25_mAd434_2 CB@25_mAd435_1 CB@25_mAd435_2 CB@25_mAd436_1 CB@25_mAd436_2 CB@25_mAd437_1 CB@25_mAd437_2 CB@25_mAd440_1 
+CB@25_mAd440_2 CB@25_mAd441_1 CB@25_mAd441_2 CB@25_mAd442_1 CB@25_mAd442_2 CB@25_mAd443_1 CB@25_mAd443_2 CB@25_mAd444_1 CB@25_mAd444_2 CB@25_mAd445_1 CB@25_mAd445_2 CB@25_mAd446_1 CB@25_mAd446_2 CB@25_mAd447_1 CB@25_mAd447_2 CB@25_mAd450_1 CB@25_mAd450_2 CB@25_mAd451_1 CB@25_mAd451_2 CB@25_mAd452_1 CB@25_mAd452_2 CB@25_mAd453_1 CB@25_mAd453_2 CB@25_mAd454_1 CB@25_mAd454_2 CB@25_mAd455_1 CB@25_mAd455_2 CB@25_mAd456_1 CB@25_mAd456_2 CB@25_mAd457_1 CB@25_mAd457_2 CB@25_mAd460_1 CB@25_mAd460_2 CB@25_mAd466_1 
+CB@25_mAd466_2 CB@25_mAd467_1 CB@25_mAd467_2 CB@25_mAd500_1 CB@25_mAd500_2 CB@25_mAd501_1 CB@25_mAd501_2 CB@25_mAd502_1 CB@25_mAd502_2 CB@25_mAd508_1 CB@25_mAd508_2 CB@25_mAd509_1 CB@25_mAd509_2 CB@25_mAd512_1 CB@25_mAd512_2 CB@25_mAd513_1 CB@25_mAd513_2 CB@25_mAd514_1 CB@25_mAd514_2 CB@25_mAd515_1 CB@25_mAd515_2 CB@25_mAd516_1 CB@25_mAd516_2 CB@25_mAd517_1 CB@25_mAd517_2 CB@25_mAd520_1 CB@25_mAd520_2 CB@25_mAd521_1 CB@25_mAd521_2 CB@25_mAd522_1 CB@25_mAd522_2 CB@25_mAd523_1 CB@25_mAd523_2 CB@25_mAd524_1 
+CB@25_mAd524_2 CB@25_mAd525_1 CB@25_mAd525_2 CB@25_mAd526_1 CB@25_mAd526_2 CB@25_mAd527_1 CB@25_mAd527_2 CB@25_mAd530_1 CB@25_mAd530_2 CB@25_mAd531_1 CB@25_mAd531_2 CB@25_mAd532_1 CB@25_mAd532_2 CB@25_mAd533_1 CB@25_mAd533_2 CB@25_mAd534_1 CB@25_mAd534_2 CB@25_mAd535_1 CB@25_mAd535_2 CB@25_mAd536_1 CB@25_mAd536_2 CB@25_mAd537_1 CB@25_mAd537_2 CB@25_mAd540_1 CB@25_mAd540_2 CB@25_mAd541_1 CB@25_mAd541_2 CB@25_mAd542_1 CB@25_mAd542_2 CB@25_mAd543_1 CB@25_mAd543_2 CB@25_mAd544_1 CB@25_mAd544_2 CB@25_mAd545_1 
+CB@25_mAd545_2 CB@25_mAd546_1 CB@25_mAd546_2 CB@25_mAd547_1 CB@25_mAd547_2 CB@25_mAd550_1 CB@25_mAd550_2 CB@25_mAd551_1 CB@25_mAd551_2 CB@25_mAd552_1 CB@25_mAd552_2 CB@25_mAd553_1 CB@25_mAd553_2 CB@25_mAd554_1 CB@25_mAd554_2 CB@25_mAd555_1 CB@25_mAd555_2 CB@25_mAd556_1 CB@25_mAd556_2 CB@25_mAd557_1 CB@25_mAd557_2 CB@25_mAd560_1 CB@25_mAd560_2 CB@25_mAd561_1 CB@25_mAd561_2 CB@25_mAd562_1 CB@25_mAd562_2 CB@25_mAd563_1 CB@25_mAd563_2 CB@25_mAd564_1 CB@25_mAd564_2 CB@25_mAd565_1 CB@25_mAd565_2 CB@25_mAd566_1 
+CB@25_mAd566_2 CB@25_mAd567_1 CB@25_mAd567_2 CB@25_mAd570_1 CB@25_mAd570_2 CB@25_mAd571_1 CB@25_mAd571_2 CB@25_mAd572_1 CB@25_mAd572_2 CB@25_mAd573_1 CB@25_mAd573_2 CB@25_mAd575_1 CB@25_mAd575_2 CB@25_mAd576_1 CB@25_mAd576_2 CB@25_mAd577_1 CB@25_mAd577_2 CB@25_mAd600_1 CB@25_mAd600_2 CB@25_mAd601_1 CB@25_mAd601_2 CB@25_mAd602_1 CB@25_mAd602_2 CB@25_mAd604_1 CB@25_mAd604_2 CB@25_mAd605_1 CB@25_mAd605_2 CB@25_mAd606_1 CB@25_mAd606_2 CB@25_mAd607_1 CB@25_mAd607_2 CB@25_mAd610_1 CB@25_mAd610_2 CB@25_mAd611_1 
+CB@25_mAd611_2 CB@25_mAd612_1 CB@25_mAd612_2 CB@25_mAd613_1 CB@25_mAd613_2 CB@25_mAd614_1 CB@25_mAd614_2 CB@25_mAd615_1 CB@25_mAd615_2 CB@25_mAd616_1 CB@25_mAd616_2 CB@25_mAd617_1 CB@25_mAd617_2 CB@25_mAd620_1 CB@25_mAd620_2 CB@25_mAd621_1 CB@25_mAd621_2 CB@25_mAd622_1 CB@25_mAd622_2 CB@25_mAd623_1 CB@25_mAd623_2 CB@25_mAd624_1 CB@25_mAd624_2 CB@25_mAd625_1 CB@25_mAd625_2 CB@25_mAd626_1 CB@25_mAd626_2 CB@25_mAd627_1 CB@25_mAd627_2 CB@25_mAd630_1 CB@25_mAd630_2 CB@25_mAd631_1 CB@25_mAd631_2 CB@25_mAd632_1 
+CB@25_mAd632_2 CB@25_mAd633_1 CB@25_mAd633_2 CB@25_mAd634_1 CB@25_mAd634_2 CB@25_mAd635_1 CB@25_mAd635_2 CB@25_mAd636_1 CB@25_mAd636_2 CB@25_mAd637_1 CB@25_mAd637_2 CB@25_mAd640_1 CB@25_mAd640_2 CB@25_mAd641_1 CB@25_mAd641_2 CB@25_mAd642_1 CB@25_mAd642_2 CB@25_mAd643_1 CB@25_mAd643_2 CB@25_mAd644_1 CB@25_mAd644_2 CB@25_mAd645_1 CB@25_mAd645_2 CB@25_mAd646_1 CB@25_mAd646_2 CB@25_mAd647_1 CB@25_mAd647_2 CB@25_mAd650_1 CB@25_mAd650_2 CB@25_mAd651_1 CB@25_mAd651_2 CB@25_mAd652_1 CB@25_mAd652_2 CB@25_mAd653_1 
+CB@25_mAd653_2 CB@25_mAd654_1 CB@25_mAd654_2 CB@25_mAd655_1 CB@25_mAd655_2 CB@25_mAd656_1 CB@25_mAd656_2 CB@25_mAd657_1 CB@25_mAd657_2 CB@25_mAd660_1 CB@25_mAd660_2 CB@25_mAd661_1 CB@25_mAd661_2 CB@25_mAd662_1 CB@25_mAd662_2 CB@25_mAd663_1 CB@25_mAd663_2 CB@25_mAd664_1 CB@25_mAd664_2 CB@25_mAd665_1 CB@25_mAd665_2 CB@25_mAd666_1 CB@25_mAd666_2 CB@25_mAd667_1 CB@25_mAd667_2 CB@25_mAd675_1 CB@25_mAd675_2 CB@25_mAd676_1 CB@25_mAd676_2 CB@25_mAd677_1 CB@25_mAd677_2 CB@25_mAd700_1 CB@25_mAd700_2 CB@25_mAd710_1 
+CB@25_mAd710_2 CB@25_mAd711_1 CB@25_mAd711_2 CB@25_mAd717_1 CB@25_mAd717_2 CB@25_mAd720_1 CB@25_mAd720_2 CB@25_mAd721_1 CB@25_mAd721_2 CB@25_mAd722_1 CB@25_mAd722_2 CB@25_mAd723_1 CB@25_mAd723_2 CB@25_mAd724_1 CB@25_mAd724_2 CB@25_mAd725_1 CB@25_mAd725_2 CB@25_mAd726_1 CB@25_mAd726_2 CB@25_mAd727_1 CB@25_mAd727_2 CB@25_mAd730_1 CB@25_mAd730_2 CB@25_mAd731_1 CB@25_mAd731_2 CB@25_mAd732_1 CB@25_mAd732_2 CB@25_mAd733_1 CB@25_mAd733_2 CB@25_mAd734_1 CB@25_mAd734_2 CB@25_mAd735_1 CB@25_mAd735_2 CB@25_mAd736_1 
+CB@25_mAd736_2 CB@25_mAd737_1 CB@25_mAd737_2 CB@25_mAd740_1 CB@25_mAd740_2 CB@25_mAd741_1 CB@25_mAd741_2 CB@25_mAd742_1 CB@25_mAd742_2 CB@25_mAd743_1 CB@25_mAd743_2 CB@25_mAd744_1 CB@25_mAd744_2 CB@25_mAd745_1 CB@25_mAd745_2 CB@25_mAd746_1 CB@25_mAd746_2 CB@25_mAd747_1 CB@25_mAd747_2 CB@25_mAd750_1 CB@25_mAd750_2 CB@25_mAd751_1 CB@25_mAd751_2 CB@25_mAd752_1 CB@25_mAd752_2 CB@25_mAd753_1 CB@25_mAd753_2 CB@25_mAd754_1 CB@25_mAd754_2 CB@25_mAd755_1 CB@25_mAd755_2 CB@25_mAd756_1 CB@25_mAd756_2 CB@25_mAd757_1 
+CB@25_mAd757_2 CB@25_mAd760_1 CB@25_mAd760_2 CB@25_mAd761_1 CB@25_mAd761_2 CB@25_mAd762_1 CB@25_mAd762_2 CB@25_mAd763_1 CB@25_mAd763_2 CB@25_mAd764_1 CB@25_mAd764_2 CB@25_mAd765_1 CB@25_mAd765_2 CB@25_mAd766_1 CB@25_mAd766_2 CB@25_mAd767_1 CB@25_mAd767_2 CB@25_mAd771_1 CB@25_mAd771_2 CB@25_mAd772_1 CB@25_mAd772_2 CB@25_mAd773_1 CB@25_mAd773_2 CB@25_mAd774_1 CB@25_mAd774_2 CB@25_mAd775_1 CB@25_mAd775_2 CB@25_mAd776_1 CB@25_mAd776_2 CB@25_mAd777_1 CB@25_mAd777_2 CB@25_X0 CB@25_X1 CB@25_X10 CB@25_X11 
+CB@25_X12 CB@25_X13 CB@25_X2 CB@25_X3 CB@25_X4 CB@25_X5 CB@25_X6 CB@25_X7 CB@25_X8 CB@25_X9 CB@25_Y1 CB@25_Y10 CB@25_Y11 CB@25_Y12 CB@25_Y2 CB@25_Y3 CB@25_Y4 CB@25_Y5 CB@25_Y6 CB@25_Y7 CB@25_Y8 CB@25_Y9 CB@25_Z1 CB@25_Z10 CB@25_Z11 CB@25_Z12 CB@25_Z2 CB@25_Z3 CB@25_Z4 CB@25_Z5 CB@25_Z6 CB@25_Z7 CB@25_Z8 CB@25_Z9 _5400TP094__CB
XCB@26 CB@26_K0 CB@26_K1 CB@26_K10 CB@26_K11 CB@26_K12 CB@26_K13 CB@26_K2 CB@26_K3 CB@26_K4 CB@26_K5 CB@26_K6 CB@26_K7 CB@26_K8 CB@26_K9 CB@26_mAd000_1 CB@26_mAd000_2 CB@26_mAd001_1 CB@26_mAd001_2 CB@26_mAd002_1 CB@26_mAd002_2 CB@26_mAd003_1 CB@26_mAd003_2 CB@26_mAd004_1 CB@26_mAd004_2 CB@26_mAd005_1 CB@26_mAd005_2 CB@26_mAd006_1 CB@26_mAd006_2 CB@26_mAd007_1 CB@26_mAd007_2 CB@26_mAd010_1 CB@26_mAd010_2 CB@26_mAd011_1 CB@26_mAd011_2 CB@26_mAd012_1 CB@26_mAd012_2 CB@26_mAd013_1 CB@26_mAd013_2 CB@26_mAd014_1 
+CB@26_mAd014_2 CB@26_mAd015_1 CB@26_mAd015_2 CB@26_mAd016_1 CB@26_mAd016_2 CB@26_mAd017_1 CB@26_mAd017_2 CB@26_mAd020_1 CB@26_mAd020_2 CB@26_mAd021_1 CB@26_mAd021_2 CB@26_mAd022_1 CB@26_mAd022_2 CB@26_mAd023_1 CB@26_mAd023_2 CB@26_mAd024_1 CB@26_mAd024_2 CB@26_mAd025_1 CB@26_mAd025_2 CB@26_mAd026_1 CB@26_mAd026_2 CB@26_mAd027_1 CB@26_mAd027_2 CB@26_mAd030_1 CB@26_mAd030_2 CB@26_mAd031_1 CB@26_mAd031_2 CB@26_mAd032_1 CB@26_mAd032_2 CB@26_mAd033_1 CB@26_mAd033_2 CB@26_mAd034_1 CB@26_mAd034_2 CB@26_mAd035_1 
+CB@26_mAd035_2 CB@26_mAd036_1 CB@26_mAd036_2 CB@26_mAd037_1 CB@26_mAd037_2 CB@26_mAd040_1 CB@26_mAd040_2 CB@26_mAd041_1 CB@26_mAd041_2 CB@26_mAd042_1 CB@26_mAd042_2 CB@26_mAd043_1 CB@26_mAd043_2 CB@26_mAd044_1 CB@26_mAd044_2 CB@26_mAd045_1 CB@26_mAd045_2 CB@26_mAd046_1 CB@26_mAd046_2 CB@26_mAd047_1 CB@26_mAd047_2 CB@26_mAd050_1 CB@26_mAd050_2 CB@26_mAd051_1 CB@26_mAd051_2 CB@26_mAd052_1 CB@26_mAd052_2 CB@26_mAd053_1 CB@26_mAd053_2 CB@26_mAd054_1 CB@26_mAd054_2 CB@26_mAd055_1 CB@26_mAd055_2 CB@26_mAd056_1 
+CB@26_mAd056_2 CB@26_mAd057_1 CB@26_mAd057_2 CB@26_mAd060_1 CB@26_mAd060_2 CB@26_mAd066_1 CB@26_mAd066_2 CB@26_mAd067_1 CB@26_mAd067_2 CB@26_mAd100_1 CB@26_mAd100_2 CB@26_mAd101_1 CB@26_mAd101_2 CB@26_mAd102_1 CB@26_mAd102_2 CB@26_mAd110_1 CB@26_mAd110_2 CB@26_mAd111_1 CB@26_mAd111_2 CB@26_mAd112_1 CB@26_mAd112_2 CB@26_mAd113_1 CB@26_mAd113_2 CB@26_mAd114_1 CB@26_mAd114_2 CB@26_mAd115_1 CB@26_mAd115_2 CB@26_mAd116_1 CB@26_mAd116_2 CB@26_mAd117_1 CB@26_mAd117_2 CB@26_mAd120_1 CB@26_mAd120_2 CB@26_mAd121_1 
+CB@26_mAd121_2 CB@26_mAd122_1 CB@26_mAd122_2 CB@26_mAd123_1 CB@26_mAd123_2 CB@26_mAd124_1 CB@26_mAd124_2 CB@26_mAd125_1 CB@26_mAd125_2 CB@26_mAd126_1 CB@26_mAd126_2 CB@26_mAd127_1 CB@26_mAd127_2 CB@26_mAd130_1 CB@26_mAd130_2 CB@26_mAd131_1 CB@26_mAd131_2 CB@26_mAd132_1 CB@26_mAd132_2 CB@26_mAd133_1 CB@26_mAd133_2 CB@26_mAd134_1 CB@26_mAd134_2 CB@26_mAd135_1 CB@26_mAd135_2 CB@26_mAd136_1 CB@26_mAd136_2 CB@26_mAd137_1 CB@26_mAd137_2 CB@26_mAd140_1 CB@26_mAd140_2 CB@26_mAd141_1 CB@26_mAd141_2 CB@26_mAd142_1 
+CB@26_mAd142_2 CB@26_mAd143_1 CB@26_mAd143_2 CB@26_mAd144_1 CB@26_mAd144_2 CB@26_mAd145_1 CB@26_mAd145_2 CB@26_mAd146_1 CB@26_mAd146_2 CB@26_mAd147_1 CB@26_mAd147_2 CB@26_mAd150_1 CB@26_mAd150_2 CB@26_mAd151_1 CB@26_mAd151_2 CB@26_mAd152_1 CB@26_mAd152_2 CB@26_mAd153_1 CB@26_mAd153_2 CB@26_mAd154_1 CB@26_mAd154_2 CB@26_mAd155_1 CB@26_mAd155_2 CB@26_mAd156_1 CB@26_mAd156_2 CB@26_mAd157_1 CB@26_mAd157_2 CB@26_mAd160_1 CB@26_mAd160_2 CB@26_mAd161_1 CB@26_mAd161_2 CB@26_mAd162_1 CB@26_mAd162_2 CB@26_mAd163_1 
+CB@26_mAd163_2 CB@26_mAd164_1 CB@26_mAd164_2 CB@26_mAd165_1 CB@26_mAd165_2 CB@26_mAd166_1 CB@26_mAd166_2 CB@26_mAd167_1 CB@26_mAd167_2 CB@26_mAd170_1 CB@26_mAd170_2 CB@26_mAd171_1 CB@26_mAd171_2 CB@26_mAd172_1 CB@26_mAd172_2 CB@26_mAd173_1 CB@26_mAd173_2 CB@26_mAd175_1 CB@26_mAd175_2 CB@26_mAd176_1 CB@26_mAd176_2 CB@26_mAd177_1 CB@26_mAd177_2 CB@26_mAd200_1 CB@26_mAd200_2 CB@26_mAd201_1 CB@26_mAd201_2 CB@26_mAd202_1 CB@26_mAd202_2 CB@26_mAd204_1 CB@26_mAd204_2 CB@26_mAd205_1 CB@26_mAd205_2 CB@26_mAd206_1 
+CB@26_mAd206_2 CB@26_mAd207_1 CB@26_mAd207_2 CB@26_mAd210_1 CB@26_mAd210_2 CB@26_mAd211_1 CB@26_mAd211_2 CB@26_mAd212_1 CB@26_mAd212_2 CB@26_mAd213_1 CB@26_mAd213_2 CB@26_mAd214_1 CB@26_mAd214_2 CB@26_mAd215_1 CB@26_mAd215_2 CB@26_mAd216_1 CB@26_mAd216_2 CB@26_mAd217_1 CB@26_mAd217_2 CB@26_mAd220_1 CB@26_mAd220_2 CB@26_mAd221_1 CB@26_mAd221_2 CB@26_mAd222_1 CB@26_mAd222_2 CB@26_mAd223_1 CB@26_mAd223_2 CB@26_mAd224_1 CB@26_mAd224_2 CB@26_mAd225_1 CB@26_mAd225_2 CB@26_mAd226_1 CB@26_mAd226_2 CB@26_mAd227_1 
+CB@26_mAd227_2 CB@26_mAd230_1 CB@26_mAd230_2 CB@26_mAd231_1 CB@26_mAd231_2 CB@26_mAd232_1 CB@26_mAd232_2 CB@26_mAd233_1 CB@26_mAd233_2 CB@26_mAd234_1 CB@26_mAd234_2 CB@26_mAd235_1 CB@26_mAd235_2 CB@26_mAd236_1 CB@26_mAd236_2 CB@26_mAd237_1 CB@26_mAd237_2 CB@26_mAd240_1 CB@26_mAd240_2 CB@26_mAd241_1 CB@26_mAd241_2 CB@26_mAd242_1 CB@26_mAd242_2 CB@26_mAd243_1 CB@26_mAd243_2 CB@26_mAd244_1 CB@26_mAd244_2 CB@26_mAd245_1 CB@26_mAd245_2 CB@26_mAd246_1 CB@26_mAd246_2 CB@26_mAd247_1 CB@26_mAd247_2 CB@26_mAd250_1 
+CB@26_mAd250_2 CB@26_mAd251_1 CB@26_mAd251_2 CB@26_mAd252_1 CB@26_mAd252_2 CB@26_mAd253_1 CB@26_mAd253_2 CB@26_mAd254_1 CB@26_mAd254_2 CB@26_mAd255_1 CB@26_mAd255_2 CB@26_mAd256_1 CB@26_mAd256_2 CB@26_mAd257_1 CB@26_mAd257_2 CB@26_mAd260_1 CB@26_mAd260_2 CB@26_mAd261_1 CB@26_mAd261_2 CB@26_mAd262_1 CB@26_mAd262_2 CB@26_mAd263_1 CB@26_mAd263_2 CB@26_mAd264_1 CB@26_mAd264_2 CB@26_mAd265_1 CB@26_mAd265_2 CB@26_mAd266_1 CB@26_mAd266_2 CB@26_mAd267_1 CB@26_mAd267_2 CB@26_mAd275_1 CB@26_mAd275_2 CB@26_mAd276_1 
+CB@26_mAd276_2 CB@26_mAd277_1 CB@26_mAd277_2 CB@26_mAd300_1 CB@26_mAd300_2 CB@26_mAd310_1 CB@26_mAd310_2 CB@26_mAd311_1 CB@26_mAd311_2 CB@26_mAd317_1 CB@26_mAd317_2 CB@26_mAd320_1 CB@26_mAd320_2 CB@26_mAd321_1 CB@26_mAd321_2 CB@26_mAd322_1 CB@26_mAd322_2 CB@26_mAd323_1 CB@26_mAd323_2 CB@26_mAd324_1 CB@26_mAd324_2 CB@26_mAd325_1 CB@26_mAd325_2 CB@26_mAd326_1 CB@26_mAd326_2 CB@26_mAd327_1 CB@26_mAd327_2 CB@26_mAd330_1 CB@26_mAd330_2 CB@26_mAd331_1 CB@26_mAd331_2 CB@26_mAd332_1 CB@26_mAd332_2 CB@26_mAd333_1 
+CB@26_mAd333_2 CB@26_mAd334_1 CB@26_mAd334_2 CB@26_mAd335_1 CB@26_mAd335_2 CB@26_mAd336_1 CB@26_mAd336_2 CB@26_mAd337_1 CB@26_mAd337_2 CB@26_mAd340_1 CB@26_mAd340_2 CB@26_mAd341_1 CB@26_mAd341_2 CB@26_mAd342_1 CB@26_mAd342_2 CB@26_mAd343_1 CB@26_mAd343_2 CB@26_mAd344_1 CB@26_mAd344_2 CB@26_mAd345_1 CB@26_mAd345_2 CB@26_mAd346_1 CB@26_mAd346_2 CB@26_mAd347_1 CB@26_mAd347_2 CB@26_mAd350_1 CB@26_mAd350_2 CB@26_mAd351_1 CB@26_mAd351_2 CB@26_mAd352_1 CB@26_mAd352_2 CB@26_mAd353_1 CB@26_mAd353_2 CB@26_mAd354_1 
+CB@26_mAd354_2 CB@26_mAd355_1 CB@26_mAd355_2 CB@26_mAd356_1 CB@26_mAd356_2 CB@26_mAd357_1 CB@26_mAd357_2 CB@26_mAd360_1 CB@26_mAd360_2 CB@26_mAd361_1 CB@26_mAd361_2 CB@26_mAd362_1 CB@26_mAd362_2 CB@26_mAd363_1 CB@26_mAd363_2 CB@26_mAd364_1 CB@26_mAd364_2 CB@26_mAd365_1 CB@26_mAd365_2 CB@26_mAd366_1 CB@26_mAd366_2 CB@26_mAd367_1 CB@26_mAd367_2 CB@26_mAd371_1 CB@26_mAd371_2 CB@26_mAd372_1 CB@26_mAd372_2 CB@26_mAd373_1 CB@26_mAd373_2 CB@26_mAd374_1 CB@26_mAd374_2 CB@26_mAd375_1 CB@26_mAd375_2 CB@26_mAd376_1 
+CB@26_mAd376_2 CB@26_mAd377_1 CB@26_mAd377_2 CB@26_mAd400_1 CB@26_mAd400_2 CB@26_mAd401_1 CB@26_mAd401_2 CB@26_mAd402_1 CB@26_mAd402_2 CB@26_mAd403_1 CB@26_mAd403_2 CB@26_mAd404_1 CB@26_mAd404_2 CB@26_mAd405_1 CB@26_mAd405_2 CB@26_mAd406_1 CB@26_mAd406_2 CB@26_mAd407_1 CB@26_mAd407_2 CB@26_mAd410_1 CB@26_mAd410_2 CB@26_mAd411_1 CB@26_mAd411_2 CB@26_mAd412_1 CB@26_mAd412_2 CB@26_mAd413_1 CB@26_mAd413_2 CB@26_mAd414_1 CB@26_mAd414_2 CB@26_mAd415_1 CB@26_mAd415_2 CB@26_mAd416_1 CB@26_mAd416_2 CB@26_mAd417_1 
+CB@26_mAd417_2 CB@26_mAd420_1 CB@26_mAd420_2 CB@26_mAd421_1 CB@26_mAd421_2 CB@26_mAd422_1 CB@26_mAd422_2 CB@26_mAd423_1 CB@26_mAd423_2 CB@26_mAd424_1 CB@26_mAd424_2 CB@26_mAd425_1 CB@26_mAd425_2 CB@26_mAd426_1 CB@26_mAd426_2 CB@26_mAd427_1 CB@26_mAd427_2 CB@26_mAd430_1 CB@26_mAd430_2 CB@26_mAd431_1 CB@26_mAd431_2 CB@26_mAd432_1 CB@26_mAd432_2 CB@26_mAd433_1 CB@26_mAd433_2 CB@26_mAd434_1 CB@26_mAd434_2 CB@26_mAd435_1 CB@26_mAd435_2 CB@26_mAd436_1 CB@26_mAd436_2 CB@26_mAd437_1 CB@26_mAd437_2 CB@26_mAd440_1 
+CB@26_mAd440_2 CB@26_mAd441_1 CB@26_mAd441_2 CB@26_mAd442_1 CB@26_mAd442_2 CB@26_mAd443_1 CB@26_mAd443_2 CB@26_mAd444_1 CB@26_mAd444_2 CB@26_mAd445_1 CB@26_mAd445_2 CB@26_mAd446_1 CB@26_mAd446_2 CB@26_mAd447_1 CB@26_mAd447_2 CB@26_mAd450_1 CB@26_mAd450_2 CB@26_mAd451_1 CB@26_mAd451_2 CB@26_mAd452_1 CB@26_mAd452_2 CB@26_mAd453_1 CB@26_mAd453_2 CB@26_mAd454_1 CB@26_mAd454_2 CB@26_mAd455_1 CB@26_mAd455_2 CB@26_mAd456_1 CB@26_mAd456_2 CB@26_mAd457_1 CB@26_mAd457_2 CB@26_mAd460_1 CB@26_mAd460_2 CB@26_mAd466_1 
+CB@26_mAd466_2 CB@26_mAd467_1 CB@26_mAd467_2 CB@26_mAd500_1 CB@26_mAd500_2 CB@26_mAd501_1 CB@26_mAd501_2 CB@26_mAd502_1 CB@26_mAd502_2 CB@26_mAd508_1 CB@26_mAd508_2 CB@26_mAd509_1 CB@26_mAd509_2 CB@26_mAd512_1 CB@26_mAd512_2 CB@26_mAd513_1 CB@26_mAd513_2 CB@26_mAd514_1 CB@26_mAd514_2 CB@26_mAd515_1 CB@26_mAd515_2 CB@26_mAd516_1 CB@26_mAd516_2 CB@26_mAd517_1 CB@26_mAd517_2 CB@26_mAd520_1 CB@26_mAd520_2 CB@26_mAd521_1 CB@26_mAd521_2 CB@26_mAd522_1 CB@26_mAd522_2 CB@26_mAd523_1 CB@26_mAd523_2 CB@26_mAd524_1 
+CB@26_mAd524_2 CB@26_mAd525_1 CB@26_mAd525_2 CB@26_mAd526_1 CB@26_mAd526_2 CB@26_mAd527_1 CB@26_mAd527_2 CB@26_mAd530_1 CB@26_mAd530_2 CB@26_mAd531_1 CB@26_mAd531_2 CB@26_mAd532_1 CB@26_mAd532_2 CB@26_mAd533_1 CB@26_mAd533_2 CB@26_mAd534_1 CB@26_mAd534_2 CB@26_mAd535_1 CB@26_mAd535_2 CB@26_mAd536_1 CB@26_mAd536_2 CB@26_mAd537_1 CB@26_mAd537_2 CB@26_mAd540_1 CB@26_mAd540_2 CB@26_mAd541_1 CB@26_mAd541_2 CB@26_mAd542_1 CB@26_mAd542_2 CB@26_mAd543_1 CB@26_mAd543_2 CB@26_mAd544_1 CB@26_mAd544_2 CB@26_mAd545_1 
+CB@26_mAd545_2 CB@26_mAd546_1 CB@26_mAd546_2 CB@26_mAd547_1 CB@26_mAd547_2 CB@26_mAd550_1 CB@26_mAd550_2 CB@26_mAd551_1 CB@26_mAd551_2 CB@26_mAd552_1 CB@26_mAd552_2 CB@26_mAd553_1 CB@26_mAd553_2 CB@26_mAd554_1 CB@26_mAd554_2 CB@26_mAd555_1 CB@26_mAd555_2 CB@26_mAd556_1 CB@26_mAd556_2 CB@26_mAd557_1 CB@26_mAd557_2 CB@26_mAd560_1 CB@26_mAd560_2 CB@26_mAd561_1 CB@26_mAd561_2 CB@26_mAd562_1 CB@26_mAd562_2 CB@26_mAd563_1 CB@26_mAd563_2 CB@26_mAd564_1 CB@26_mAd564_2 CB@26_mAd565_1 CB@26_mAd565_2 CB@26_mAd566_1 
+CB@26_mAd566_2 CB@26_mAd567_1 CB@26_mAd567_2 CB@26_mAd570_1 CB@26_mAd570_2 CB@26_mAd571_1 CB@26_mAd571_2 CB@26_mAd572_1 CB@26_mAd572_2 CB@26_mAd573_1 CB@26_mAd573_2 CB@26_mAd575_1 CB@26_mAd575_2 CB@26_mAd576_1 CB@26_mAd576_2 CB@26_mAd577_1 CB@26_mAd577_2 CB@26_mAd600_1 CB@26_mAd600_2 CB@26_mAd601_1 CB@26_mAd601_2 CB@26_mAd602_1 CB@26_mAd602_2 CB@26_mAd604_1 CB@26_mAd604_2 CB@26_mAd605_1 CB@26_mAd605_2 CB@26_mAd606_1 CB@26_mAd606_2 CB@26_mAd607_1 CB@26_mAd607_2 CB@26_mAd610_1 CB@26_mAd610_2 CB@26_mAd611_1 
+CB@26_mAd611_2 CB@26_mAd612_1 CB@26_mAd612_2 CB@26_mAd613_1 CB@26_mAd613_2 CB@26_mAd614_1 CB@26_mAd614_2 CB@26_mAd615_1 CB@26_mAd615_2 CB@26_mAd616_1 CB@26_mAd616_2 CB@26_mAd617_1 CB@26_mAd617_2 CB@26_mAd620_1 CB@26_mAd620_2 CB@26_mAd621_1 CB@26_mAd621_2 CB@26_mAd622_1 CB@26_mAd622_2 CB@26_mAd623_1 CB@26_mAd623_2 CB@26_mAd624_1 CB@26_mAd624_2 CB@26_mAd625_1 CB@26_mAd625_2 CB@26_mAd626_1 CB@26_mAd626_2 CB@26_mAd627_1 CB@26_mAd627_2 CB@26_mAd630_1 CB@26_mAd630_2 CB@26_mAd631_1 CB@26_mAd631_2 CB@26_mAd632_1 
+CB@26_mAd632_2 CB@26_mAd633_1 CB@26_mAd633_2 CB@26_mAd634_1 CB@26_mAd634_2 CB@26_mAd635_1 CB@26_mAd635_2 CB@26_mAd636_1 CB@26_mAd636_2 CB@26_mAd637_1 CB@26_mAd637_2 CB@26_mAd640_1 CB@26_mAd640_2 CB@26_mAd641_1 CB@26_mAd641_2 CB@26_mAd642_1 CB@26_mAd642_2 CB@26_mAd643_1 CB@26_mAd643_2 CB@26_mAd644_1 CB@26_mAd644_2 CB@26_mAd645_1 CB@26_mAd645_2 CB@26_mAd646_1 CB@26_mAd646_2 CB@26_mAd647_1 CB@26_mAd647_2 CB@26_mAd650_1 CB@26_mAd650_2 CB@26_mAd651_1 CB@26_mAd651_2 CB@26_mAd652_1 CB@26_mAd652_2 CB@26_mAd653_1 
+CB@26_mAd653_2 CB@26_mAd654_1 CB@26_mAd654_2 CB@26_mAd655_1 CB@26_mAd655_2 CB@26_mAd656_1 CB@26_mAd656_2 CB@26_mAd657_1 CB@26_mAd657_2 CB@26_mAd660_1 CB@26_mAd660_2 CB@26_mAd661_1 CB@26_mAd661_2 CB@26_mAd662_1 CB@26_mAd662_2 CB@26_mAd663_1 CB@26_mAd663_2 CB@26_mAd664_1 CB@26_mAd664_2 CB@26_mAd665_1 CB@26_mAd665_2 CB@26_mAd666_1 CB@26_mAd666_2 CB@26_mAd667_1 CB@26_mAd667_2 CB@26_mAd675_1 CB@26_mAd675_2 CB@26_mAd676_1 CB@26_mAd676_2 CB@26_mAd677_1 CB@26_mAd677_2 CB@26_mAd700_1 CB@26_mAd700_2 CB@26_mAd710_1 
+CB@26_mAd710_2 CB@26_mAd711_1 CB@26_mAd711_2 CB@26_mAd717_1 CB@26_mAd717_2 CB@26_mAd720_1 CB@26_mAd720_2 CB@26_mAd721_1 CB@26_mAd721_2 CB@26_mAd722_1 CB@26_mAd722_2 CB@26_mAd723_1 CB@26_mAd723_2 CB@26_mAd724_1 CB@26_mAd724_2 CB@26_mAd725_1 CB@26_mAd725_2 CB@26_mAd726_1 CB@26_mAd726_2 CB@26_mAd727_1 CB@26_mAd727_2 CB@26_mAd730_1 CB@26_mAd730_2 CB@26_mAd731_1 CB@26_mAd731_2 CB@26_mAd732_1 CB@26_mAd732_2 CB@26_mAd733_1 CB@26_mAd733_2 CB@26_mAd734_1 CB@26_mAd734_2 CB@26_mAd735_1 CB@26_mAd735_2 CB@26_mAd736_1 
+CB@26_mAd736_2 CB@26_mAd737_1 CB@26_mAd737_2 CB@26_mAd740_1 CB@26_mAd740_2 CB@26_mAd741_1 CB@26_mAd741_2 CB@26_mAd742_1 CB@26_mAd742_2 CB@26_mAd743_1 CB@26_mAd743_2 CB@26_mAd744_1 CB@26_mAd744_2 CB@26_mAd745_1 CB@26_mAd745_2 CB@26_mAd746_1 CB@26_mAd746_2 CB@26_mAd747_1 CB@26_mAd747_2 CB@26_mAd750_1 CB@26_mAd750_2 CB@26_mAd751_1 CB@26_mAd751_2 CB@26_mAd752_1 CB@26_mAd752_2 CB@26_mAd753_1 CB@26_mAd753_2 CB@26_mAd754_1 CB@26_mAd754_2 CB@26_mAd755_1 CB@26_mAd755_2 CB@26_mAd756_1 CB@26_mAd756_2 CB@26_mAd757_1 
+CB@26_mAd757_2 CB@26_mAd760_1 CB@26_mAd760_2 CB@26_mAd761_1 CB@26_mAd761_2 CB@26_mAd762_1 CB@26_mAd762_2 CB@26_mAd763_1 CB@26_mAd763_2 CB@26_mAd764_1 CB@26_mAd764_2 CB@26_mAd765_1 CB@26_mAd765_2 CB@26_mAd766_1 CB@26_mAd766_2 CB@26_mAd767_1 CB@26_mAd767_2 CB@26_mAd771_1 CB@26_mAd771_2 CB@26_mAd772_1 CB@26_mAd772_2 CB@26_mAd773_1 CB@26_mAd773_2 CB@26_mAd774_1 CB@26_mAd774_2 CB@26_mAd775_1 CB@26_mAd775_2 CB@26_mAd776_1 CB@26_mAd776_2 CB@26_mAd777_1 CB@26_mAd777_2 CB@26_X0 CB@26_X1 CB@26_X10 CB@26_X11 
+CB@26_X12 CB@26_X13 CB@26_X2 CB@26_X3 CB@26_X4 CB@26_X5 CB@26_X6 CB@26_X7 CB@26_X8 CB@26_X9 CB@26_Y1 CB@26_Y10 CB@26_Y11 CB@26_Y12 CB@26_Y2 CB@26_Y3 CB@26_Y4 CB@26_Y5 CB@26_Y6 CB@26_Y7 CB@26_Y8 CB@26_Y9 CB@26_Z1 CB@26_Z10 CB@26_Z11 CB@26_Z12 CB@26_Z2 CB@26_Z3 CB@26_Z4 CB@26_Z5 CB@26_Z6 CB@26_Z7 CB@26_Z8 CB@26_Z9 _5400TP094__CB
XCB@27 CB@27_K0 CB@27_K1 CB@27_K10 CB@27_K11 CB@27_K12 CB@27_K13 CB@27_K2 CB@27_K3 CB@27_K4 CB@27_K5 CB@27_K6 CB@27_K7 CB@27_K8 CB@27_K9 CB@27_mAd000_1 CB@27_mAd000_2 CB@27_mAd001_1 CB@27_mAd001_2 CB@27_mAd002_1 CB@27_mAd002_2 CB@27_mAd003_1 CB@27_mAd003_2 CB@27_mAd004_1 CB@27_mAd004_2 CB@27_mAd005_1 CB@27_mAd005_2 CB@27_mAd006_1 CB@27_mAd006_2 CB@27_mAd007_1 CB@27_mAd007_2 CB@27_mAd010_1 CB@27_mAd010_2 CB@27_mAd011_1 CB@27_mAd011_2 CB@27_mAd012_1 CB@27_mAd012_2 CB@27_mAd013_1 CB@27_mAd013_2 CB@27_mAd014_1 
+CB@27_mAd014_2 CB@27_mAd015_1 CB@27_mAd015_2 CB@27_mAd016_1 CB@27_mAd016_2 CB@27_mAd017_1 CB@27_mAd017_2 CB@27_mAd020_1 CB@27_mAd020_2 CB@27_mAd021_1 CB@27_mAd021_2 CB@27_mAd022_1 CB@27_mAd022_2 CB@27_mAd023_1 CB@27_mAd023_2 CB@27_mAd024_1 CB@27_mAd024_2 CB@27_mAd025_1 CB@27_mAd025_2 CB@27_mAd026_1 CB@27_mAd026_2 CB@27_mAd027_1 CB@27_mAd027_2 CB@27_mAd030_1 CB@27_mAd030_2 CB@27_mAd031_1 CB@27_mAd031_2 CB@27_mAd032_1 CB@27_mAd032_2 CB@27_mAd033_1 CB@27_mAd033_2 CB@27_mAd034_1 CB@27_mAd034_2 CB@27_mAd035_1 
+CB@27_mAd035_2 CB@27_mAd036_1 CB@27_mAd036_2 CB@27_mAd037_1 CB@27_mAd037_2 CB@27_mAd040_1 CB@27_mAd040_2 CB@27_mAd041_1 CB@27_mAd041_2 CB@27_mAd042_1 CB@27_mAd042_2 CB@27_mAd043_1 CB@27_mAd043_2 CB@27_mAd044_1 CB@27_mAd044_2 CB@27_mAd045_1 CB@27_mAd045_2 CB@27_mAd046_1 CB@27_mAd046_2 CB@27_mAd047_1 CB@27_mAd047_2 CB@27_mAd050_1 CB@27_mAd050_2 CB@27_mAd051_1 CB@27_mAd051_2 CB@27_mAd052_1 CB@27_mAd052_2 CB@27_mAd053_1 CB@27_mAd053_2 CB@27_mAd054_1 CB@27_mAd054_2 CB@27_mAd055_1 CB@27_mAd055_2 CB@27_mAd056_1 
+CB@27_mAd056_2 CB@27_mAd057_1 CB@27_mAd057_2 CB@27_mAd060_1 CB@27_mAd060_2 CB@27_mAd066_1 CB@27_mAd066_2 CB@27_mAd067_1 CB@27_mAd067_2 CB@27_mAd100_1 CB@27_mAd100_2 CB@27_mAd101_1 CB@27_mAd101_2 CB@27_mAd102_1 CB@27_mAd102_2 CB@27_mAd110_1 CB@27_mAd110_2 CB@27_mAd111_1 CB@27_mAd111_2 CB@27_mAd112_1 CB@27_mAd112_2 CB@27_mAd113_1 CB@27_mAd113_2 CB@27_mAd114_1 CB@27_mAd114_2 CB@27_mAd115_1 CB@27_mAd115_2 CB@27_mAd116_1 CB@27_mAd116_2 CB@27_mAd117_1 CB@27_mAd117_2 CB@27_mAd120_1 CB@27_mAd120_2 CB@27_mAd121_1 
+CB@27_mAd121_2 CB@27_mAd122_1 CB@27_mAd122_2 CB@27_mAd123_1 CB@27_mAd123_2 CB@27_mAd124_1 CB@27_mAd124_2 CB@27_mAd125_1 CB@27_mAd125_2 CB@27_mAd126_1 CB@27_mAd126_2 CB@27_mAd127_1 CB@27_mAd127_2 CB@27_mAd130_1 CB@27_mAd130_2 CB@27_mAd131_1 CB@27_mAd131_2 CB@27_mAd132_1 CB@27_mAd132_2 CB@27_mAd133_1 CB@27_mAd133_2 CB@27_mAd134_1 CB@27_mAd134_2 CB@27_mAd135_1 CB@27_mAd135_2 CB@27_mAd136_1 CB@27_mAd136_2 CB@27_mAd137_1 CB@27_mAd137_2 CB@27_mAd140_1 CB@27_mAd140_2 CB@27_mAd141_1 CB@27_mAd141_2 CB@27_mAd142_1 
+CB@27_mAd142_2 CB@27_mAd143_1 CB@27_mAd143_2 CB@27_mAd144_1 CB@27_mAd144_2 CB@27_mAd145_1 CB@27_mAd145_2 CB@27_mAd146_1 CB@27_mAd146_2 CB@27_mAd147_1 CB@27_mAd147_2 CB@27_mAd150_1 CB@27_mAd150_2 CB@27_mAd151_1 CB@27_mAd151_2 CB@27_mAd152_1 CB@27_mAd152_2 CB@27_mAd153_1 CB@27_mAd153_2 CB@27_mAd154_1 CB@27_mAd154_2 CB@27_mAd155_1 CB@27_mAd155_2 CB@27_mAd156_1 CB@27_mAd156_2 CB@27_mAd157_1 CB@27_mAd157_2 CB@27_mAd160_1 CB@27_mAd160_2 CB@27_mAd161_1 CB@27_mAd161_2 CB@27_mAd162_1 CB@27_mAd162_2 CB@27_mAd163_1 
+CB@27_mAd163_2 CB@27_mAd164_1 CB@27_mAd164_2 CB@27_mAd165_1 CB@27_mAd165_2 CB@27_mAd166_1 CB@27_mAd166_2 CB@27_mAd167_1 CB@27_mAd167_2 CB@27_mAd170_1 CB@27_mAd170_2 CB@27_mAd171_1 CB@27_mAd171_2 CB@27_mAd172_1 CB@27_mAd172_2 CB@27_mAd173_1 CB@27_mAd173_2 CB@27_mAd175_1 CB@27_mAd175_2 CB@27_mAd176_1 CB@27_mAd176_2 CB@27_mAd177_1 CB@27_mAd177_2 CB@27_mAd200_1 CB@27_mAd200_2 CB@27_mAd201_1 CB@27_mAd201_2 CB@27_mAd202_1 CB@27_mAd202_2 CB@27_mAd204_1 CB@27_mAd204_2 CB@27_mAd205_1 CB@27_mAd205_2 CB@27_mAd206_1 
+CB@27_mAd206_2 CB@27_mAd207_1 CB@27_mAd207_2 CB@27_mAd210_1 CB@27_mAd210_2 CB@27_mAd211_1 CB@27_mAd211_2 CB@27_mAd212_1 CB@27_mAd212_2 CB@27_mAd213_1 CB@27_mAd213_2 CB@27_mAd214_1 CB@27_mAd214_2 CB@27_mAd215_1 CB@27_mAd215_2 CB@27_mAd216_1 CB@27_mAd216_2 CB@27_mAd217_1 CB@27_mAd217_2 CB@27_mAd220_1 CB@27_mAd220_2 CB@27_mAd221_1 CB@27_mAd221_2 CB@27_mAd222_1 CB@27_mAd222_2 CB@27_mAd223_1 CB@27_mAd223_2 CB@27_mAd224_1 CB@27_mAd224_2 CB@27_mAd225_1 CB@27_mAd225_2 CB@27_mAd226_1 CB@27_mAd226_2 CB@27_mAd227_1 
+CB@27_mAd227_2 CB@27_mAd230_1 CB@27_mAd230_2 CB@27_mAd231_1 CB@27_mAd231_2 CB@27_mAd232_1 CB@27_mAd232_2 CB@27_mAd233_1 CB@27_mAd233_2 CB@27_mAd234_1 CB@27_mAd234_2 CB@27_mAd235_1 CB@27_mAd235_2 CB@27_mAd236_1 CB@27_mAd236_2 CB@27_mAd237_1 CB@27_mAd237_2 CB@27_mAd240_1 CB@27_mAd240_2 CB@27_mAd241_1 CB@27_mAd241_2 CB@27_mAd242_1 CB@27_mAd242_2 CB@27_mAd243_1 CB@27_mAd243_2 CB@27_mAd244_1 CB@27_mAd244_2 CB@27_mAd245_1 CB@27_mAd245_2 CB@27_mAd246_1 CB@27_mAd246_2 CB@27_mAd247_1 CB@27_mAd247_2 CB@27_mAd250_1 
+CB@27_mAd250_2 CB@27_mAd251_1 CB@27_mAd251_2 CB@27_mAd252_1 CB@27_mAd252_2 CB@27_mAd253_1 CB@27_mAd253_2 CB@27_mAd254_1 CB@27_mAd254_2 CB@27_mAd255_1 CB@27_mAd255_2 CB@27_mAd256_1 CB@27_mAd256_2 CB@27_mAd257_1 CB@27_mAd257_2 CB@27_mAd260_1 CB@27_mAd260_2 CB@27_mAd261_1 CB@27_mAd261_2 CB@27_mAd262_1 CB@27_mAd262_2 CB@27_mAd263_1 CB@27_mAd263_2 CB@27_mAd264_1 CB@27_mAd264_2 CB@27_mAd265_1 CB@27_mAd265_2 CB@27_mAd266_1 CB@27_mAd266_2 CB@27_mAd267_1 CB@27_mAd267_2 CB@27_mAd275_1 CB@27_mAd275_2 CB@27_mAd276_1 
+CB@27_mAd276_2 CB@27_mAd277_1 CB@27_mAd277_2 CB@27_mAd300_1 CB@27_mAd300_2 CB@27_mAd310_1 CB@27_mAd310_2 CB@27_mAd311_1 CB@27_mAd311_2 CB@27_mAd317_1 CB@27_mAd317_2 CB@27_mAd320_1 CB@27_mAd320_2 CB@27_mAd321_1 CB@27_mAd321_2 CB@27_mAd322_1 CB@27_mAd322_2 CB@27_mAd323_1 CB@27_mAd323_2 CB@27_mAd324_1 CB@27_mAd324_2 CB@27_mAd325_1 CB@27_mAd325_2 CB@27_mAd326_1 CB@27_mAd326_2 CB@27_mAd327_1 CB@27_mAd327_2 CB@27_mAd330_1 CB@27_mAd330_2 CB@27_mAd331_1 CB@27_mAd331_2 CB@27_mAd332_1 CB@27_mAd332_2 CB@27_mAd333_1 
+CB@27_mAd333_2 CB@27_mAd334_1 CB@27_mAd334_2 CB@27_mAd335_1 CB@27_mAd335_2 CB@27_mAd336_1 CB@27_mAd336_2 CB@27_mAd337_1 CB@27_mAd337_2 CB@27_mAd340_1 CB@27_mAd340_2 CB@27_mAd341_1 CB@27_mAd341_2 CB@27_mAd342_1 CB@27_mAd342_2 CB@27_mAd343_1 CB@27_mAd343_2 CB@27_mAd344_1 CB@27_mAd344_2 CB@27_mAd345_1 CB@27_mAd345_2 CB@27_mAd346_1 CB@27_mAd346_2 CB@27_mAd347_1 CB@27_mAd347_2 CB@27_mAd350_1 CB@27_mAd350_2 CB@27_mAd351_1 CB@27_mAd351_2 CB@27_mAd352_1 CB@27_mAd352_2 CB@27_mAd353_1 CB@27_mAd353_2 CB@27_mAd354_1 
+CB@27_mAd354_2 CB@27_mAd355_1 CB@27_mAd355_2 CB@27_mAd356_1 CB@27_mAd356_2 CB@27_mAd357_1 CB@27_mAd357_2 CB@27_mAd360_1 CB@27_mAd360_2 CB@27_mAd361_1 CB@27_mAd361_2 CB@27_mAd362_1 CB@27_mAd362_2 CB@27_mAd363_1 CB@27_mAd363_2 CB@27_mAd364_1 CB@27_mAd364_2 CB@27_mAd365_1 CB@27_mAd365_2 CB@27_mAd366_1 CB@27_mAd366_2 CB@27_mAd367_1 CB@27_mAd367_2 CB@27_mAd371_1 CB@27_mAd371_2 CB@27_mAd372_1 CB@27_mAd372_2 CB@27_mAd373_1 CB@27_mAd373_2 CB@27_mAd374_1 CB@27_mAd374_2 CB@27_mAd375_1 CB@27_mAd375_2 CB@27_mAd376_1 
+CB@27_mAd376_2 CB@27_mAd377_1 CB@27_mAd377_2 CB@27_mAd400_1 CB@27_mAd400_2 CB@27_mAd401_1 CB@27_mAd401_2 CB@27_mAd402_1 CB@27_mAd402_2 CB@27_mAd403_1 CB@27_mAd403_2 CB@27_mAd404_1 CB@27_mAd404_2 CB@27_mAd405_1 CB@27_mAd405_2 CB@27_mAd406_1 CB@27_mAd406_2 CB@27_mAd407_1 CB@27_mAd407_2 CB@27_mAd410_1 CB@27_mAd410_2 CB@27_mAd411_1 CB@27_mAd411_2 CB@27_mAd412_1 CB@27_mAd412_2 CB@27_mAd413_1 CB@27_mAd413_2 CB@27_mAd414_1 CB@27_mAd414_2 CB@27_mAd415_1 CB@27_mAd415_2 CB@27_mAd416_1 CB@27_mAd416_2 CB@27_mAd417_1 
+CB@27_mAd417_2 CB@27_mAd420_1 CB@27_mAd420_2 CB@27_mAd421_1 CB@27_mAd421_2 CB@27_mAd422_1 CB@27_mAd422_2 CB@27_mAd423_1 CB@27_mAd423_2 CB@27_mAd424_1 CB@27_mAd424_2 CB@27_mAd425_1 CB@27_mAd425_2 CB@27_mAd426_1 CB@27_mAd426_2 CB@27_mAd427_1 CB@27_mAd427_2 CB@27_mAd430_1 CB@27_mAd430_2 CB@27_mAd431_1 CB@27_mAd431_2 CB@27_mAd432_1 CB@27_mAd432_2 CB@27_mAd433_1 CB@27_mAd433_2 CB@27_mAd434_1 CB@27_mAd434_2 CB@27_mAd435_1 CB@27_mAd435_2 CB@27_mAd436_1 CB@27_mAd436_2 CB@27_mAd437_1 CB@27_mAd437_2 CB@27_mAd440_1 
+CB@27_mAd440_2 CB@27_mAd441_1 CB@27_mAd441_2 CB@27_mAd442_1 CB@27_mAd442_2 CB@27_mAd443_1 CB@27_mAd443_2 CB@27_mAd444_1 CB@27_mAd444_2 CB@27_mAd445_1 CB@27_mAd445_2 CB@27_mAd446_1 CB@27_mAd446_2 CB@27_mAd447_1 CB@27_mAd447_2 CB@27_mAd450_1 CB@27_mAd450_2 CB@27_mAd451_1 CB@27_mAd451_2 CB@27_mAd452_1 CB@27_mAd452_2 CB@27_mAd453_1 CB@27_mAd453_2 CB@27_mAd454_1 CB@27_mAd454_2 CB@27_mAd455_1 CB@27_mAd455_2 CB@27_mAd456_1 CB@27_mAd456_2 CB@27_mAd457_1 CB@27_mAd457_2 CB@27_mAd460_1 CB@27_mAd460_2 CB@27_mAd466_1 
+CB@27_mAd466_2 CB@27_mAd467_1 CB@27_mAd467_2 CB@27_mAd500_1 CB@27_mAd500_2 CB@27_mAd501_1 CB@27_mAd501_2 CB@27_mAd502_1 CB@27_mAd502_2 CB@27_mAd508_1 CB@27_mAd508_2 CB@27_mAd509_1 CB@27_mAd509_2 CB@27_mAd512_1 CB@27_mAd512_2 CB@27_mAd513_1 CB@27_mAd513_2 CB@27_mAd514_1 CB@27_mAd514_2 CB@27_mAd515_1 CB@27_mAd515_2 CB@27_mAd516_1 CB@27_mAd516_2 CB@27_mAd517_1 CB@27_mAd517_2 CB@27_mAd520_1 CB@27_mAd520_2 CB@27_mAd521_1 CB@27_mAd521_2 CB@27_mAd522_1 CB@27_mAd522_2 CB@27_mAd523_1 CB@27_mAd523_2 CB@27_mAd524_1 
+CB@27_mAd524_2 CB@27_mAd525_1 CB@27_mAd525_2 CB@27_mAd526_1 CB@27_mAd526_2 CB@27_mAd527_1 CB@27_mAd527_2 CB@27_mAd530_1 CB@27_mAd530_2 CB@27_mAd531_1 CB@27_mAd531_2 CB@27_mAd532_1 CB@27_mAd532_2 CB@27_mAd533_1 CB@27_mAd533_2 CB@27_mAd534_1 CB@27_mAd534_2 CB@27_mAd535_1 CB@27_mAd535_2 CB@27_mAd536_1 CB@27_mAd536_2 CB@27_mAd537_1 CB@27_mAd537_2 CB@27_mAd540_1 CB@27_mAd540_2 CB@27_mAd541_1 CB@27_mAd541_2 CB@27_mAd542_1 CB@27_mAd542_2 CB@27_mAd543_1 CB@27_mAd543_2 CB@27_mAd544_1 CB@27_mAd544_2 CB@27_mAd545_1 
+CB@27_mAd545_2 CB@27_mAd546_1 CB@27_mAd546_2 CB@27_mAd547_1 CB@27_mAd547_2 CB@27_mAd550_1 CB@27_mAd550_2 CB@27_mAd551_1 CB@27_mAd551_2 CB@27_mAd552_1 CB@27_mAd552_2 CB@27_mAd553_1 CB@27_mAd553_2 CB@27_mAd554_1 CB@27_mAd554_2 CB@27_mAd555_1 CB@27_mAd555_2 CB@27_mAd556_1 CB@27_mAd556_2 CB@27_mAd557_1 CB@27_mAd557_2 CB@27_mAd560_1 CB@27_mAd560_2 CB@27_mAd561_1 CB@27_mAd561_2 CB@27_mAd562_1 CB@27_mAd562_2 CB@27_mAd563_1 CB@27_mAd563_2 CB@27_mAd564_1 CB@27_mAd564_2 CB@27_mAd565_1 CB@27_mAd565_2 CB@27_mAd566_1 
+CB@27_mAd566_2 CB@27_mAd567_1 CB@27_mAd567_2 CB@27_mAd570_1 CB@27_mAd570_2 CB@27_mAd571_1 CB@27_mAd571_2 CB@27_mAd572_1 CB@27_mAd572_2 CB@27_mAd573_1 CB@27_mAd573_2 CB@27_mAd575_1 CB@27_mAd575_2 CB@27_mAd576_1 CB@27_mAd576_2 CB@27_mAd577_1 CB@27_mAd577_2 CB@27_mAd600_1 CB@27_mAd600_2 CB@27_mAd601_1 CB@27_mAd601_2 CB@27_mAd602_1 CB@27_mAd602_2 CB@27_mAd604_1 CB@27_mAd604_2 CB@27_mAd605_1 CB@27_mAd605_2 CB@27_mAd606_1 CB@27_mAd606_2 CB@27_mAd607_1 CB@27_mAd607_2 CB@27_mAd610_1 CB@27_mAd610_2 CB@27_mAd611_1 
+CB@27_mAd611_2 CB@27_mAd612_1 CB@27_mAd612_2 CB@27_mAd613_1 CB@27_mAd613_2 CB@27_mAd614_1 CB@27_mAd614_2 CB@27_mAd615_1 CB@27_mAd615_2 CB@27_mAd616_1 CB@27_mAd616_2 CB@27_mAd617_1 CB@27_mAd617_2 CB@27_mAd620_1 CB@27_mAd620_2 CB@27_mAd621_1 CB@27_mAd621_2 CB@27_mAd622_1 CB@27_mAd622_2 CB@27_mAd623_1 CB@27_mAd623_2 CB@27_mAd624_1 CB@27_mAd624_2 CB@27_mAd625_1 CB@27_mAd625_2 CB@27_mAd626_1 CB@27_mAd626_2 CB@27_mAd627_1 CB@27_mAd627_2 CB@27_mAd630_1 CB@27_mAd630_2 CB@27_mAd631_1 CB@27_mAd631_2 CB@27_mAd632_1 
+CB@27_mAd632_2 CB@27_mAd633_1 CB@27_mAd633_2 CB@27_mAd634_1 CB@27_mAd634_2 CB@27_mAd635_1 CB@27_mAd635_2 CB@27_mAd636_1 CB@27_mAd636_2 CB@27_mAd637_1 CB@27_mAd637_2 CB@27_mAd640_1 CB@27_mAd640_2 CB@27_mAd641_1 CB@27_mAd641_2 CB@27_mAd642_1 CB@27_mAd642_2 CB@27_mAd643_1 CB@27_mAd643_2 CB@27_mAd644_1 CB@27_mAd644_2 CB@27_mAd645_1 CB@27_mAd645_2 CB@27_mAd646_1 CB@27_mAd646_2 CB@27_mAd647_1 CB@27_mAd647_2 CB@27_mAd650_1 CB@27_mAd650_2 CB@27_mAd651_1 CB@27_mAd651_2 CB@27_mAd652_1 CB@27_mAd652_2 CB@27_mAd653_1 
+CB@27_mAd653_2 CB@27_mAd654_1 CB@27_mAd654_2 CB@27_mAd655_1 CB@27_mAd655_2 CB@27_mAd656_1 CB@27_mAd656_2 CB@27_mAd657_1 CB@27_mAd657_2 CB@27_mAd660_1 CB@27_mAd660_2 CB@27_mAd661_1 CB@27_mAd661_2 CB@27_mAd662_1 CB@27_mAd662_2 CB@27_mAd663_1 CB@27_mAd663_2 CB@27_mAd664_1 CB@27_mAd664_2 CB@27_mAd665_1 CB@27_mAd665_2 CB@27_mAd666_1 CB@27_mAd666_2 CB@27_mAd667_1 CB@27_mAd667_2 CB@27_mAd675_1 CB@27_mAd675_2 CB@27_mAd676_1 CB@27_mAd676_2 CB@27_mAd677_1 CB@27_mAd677_2 CB@27_mAd700_1 CB@27_mAd700_2 CB@27_mAd710_1 
+CB@27_mAd710_2 CB@27_mAd711_1 CB@27_mAd711_2 CB@27_mAd717_1 CB@27_mAd717_2 CB@27_mAd720_1 CB@27_mAd720_2 CB@27_mAd721_1 CB@27_mAd721_2 CB@27_mAd722_1 CB@27_mAd722_2 CB@27_mAd723_1 CB@27_mAd723_2 CB@27_mAd724_1 CB@27_mAd724_2 CB@27_mAd725_1 CB@27_mAd725_2 CB@27_mAd726_1 CB@27_mAd726_2 CB@27_mAd727_1 CB@27_mAd727_2 CB@27_mAd730_1 CB@27_mAd730_2 CB@27_mAd731_1 CB@27_mAd731_2 CB@27_mAd732_1 CB@27_mAd732_2 CB@27_mAd733_1 CB@27_mAd733_2 CB@27_mAd734_1 CB@27_mAd734_2 CB@27_mAd735_1 CB@27_mAd735_2 CB@27_mAd736_1 
+CB@27_mAd736_2 CB@27_mAd737_1 CB@27_mAd737_2 CB@27_mAd740_1 CB@27_mAd740_2 CB@27_mAd741_1 CB@27_mAd741_2 CB@27_mAd742_1 CB@27_mAd742_2 CB@27_mAd743_1 CB@27_mAd743_2 CB@27_mAd744_1 CB@27_mAd744_2 CB@27_mAd745_1 CB@27_mAd745_2 CB@27_mAd746_1 CB@27_mAd746_2 CB@27_mAd747_1 CB@27_mAd747_2 CB@27_mAd750_1 CB@27_mAd750_2 CB@27_mAd751_1 CB@27_mAd751_2 CB@27_mAd752_1 CB@27_mAd752_2 CB@27_mAd753_1 CB@27_mAd753_2 CB@27_mAd754_1 CB@27_mAd754_2 CB@27_mAd755_1 CB@27_mAd755_2 CB@27_mAd756_1 CB@27_mAd756_2 CB@27_mAd757_1 
+CB@27_mAd757_2 CB@27_mAd760_1 CB@27_mAd760_2 CB@27_mAd761_1 CB@27_mAd761_2 CB@27_mAd762_1 CB@27_mAd762_2 CB@27_mAd763_1 CB@27_mAd763_2 CB@27_mAd764_1 CB@27_mAd764_2 CB@27_mAd765_1 CB@27_mAd765_2 CB@27_mAd766_1 CB@27_mAd766_2 CB@27_mAd767_1 CB@27_mAd767_2 CB@27_mAd771_1 CB@27_mAd771_2 CB@27_mAd772_1 CB@27_mAd772_2 CB@27_mAd773_1 CB@27_mAd773_2 CB@27_mAd774_1 CB@27_mAd774_2 CB@27_mAd775_1 CB@27_mAd775_2 CB@27_mAd776_1 CB@27_mAd776_2 CB@27_mAd777_1 CB@27_mAd777_2 CB@27_X0 CB@27_X1 CB@27_X10 CB@27_X11 
+CB@27_X12 CB@27_X13 CB@27_X2 CB@27_X3 CB@27_X4 CB@27_X5 CB@27_X6 CB@27_X7 CB@27_X8 CB@27_X9 CB@27_Y1 CB@27_Y10 CB@27_Y11 CB@27_Y12 CB@27_Y2 CB@27_Y3 CB@27_Y4 CB@27_Y5 CB@27_Y6 CB@27_Y7 CB@27_Y8 CB@27_Y9 CB@27_Z1 CB@27_Z10 CB@27_Z11 CB@27_Z12 CB@27_Z2 CB@27_Z3 CB@27_Z4 CB@27_Z5 CB@27_Z6 CB@27_Z7 CB@27_Z8 CB@27_Z9 _5400TP094__CB
XCB@28 CB@28_K0 CB@28_K1 CB@28_K10 CB@28_K11 CB@28_K12 CB@28_K13 CB@28_K2 CB@28_K3 CB@28_K4 CB@28_K5 CB@28_K6 CB@28_K7 CB@28_K8 CB@28_K9 CB@28_mAd000_1 CB@28_mAd000_2 CB@28_mAd001_1 CB@28_mAd001_2 CB@28_mAd002_1 CB@28_mAd002_2 CB@28_mAd003_1 CB@28_mAd003_2 CB@28_mAd004_1 CB@28_mAd004_2 CB@28_mAd005_1 CB@28_mAd005_2 CB@28_mAd006_1 CB@28_mAd006_2 CB@28_mAd007_1 CB@28_mAd007_2 CB@28_mAd010_1 CB@28_mAd010_2 CB@28_mAd011_1 CB@28_mAd011_2 CB@28_mAd012_1 CB@28_mAd012_2 CB@28_mAd013_1 CB@28_mAd013_2 CB@28_mAd014_1 
+CB@28_mAd014_2 CB@28_mAd015_1 CB@28_mAd015_2 CB@28_mAd016_1 CB@28_mAd016_2 CB@28_mAd017_1 CB@28_mAd017_2 CB@28_mAd020_1 CB@28_mAd020_2 CB@28_mAd021_1 CB@28_mAd021_2 CB@28_mAd022_1 CB@28_mAd022_2 CB@28_mAd023_1 CB@28_mAd023_2 CB@28_mAd024_1 CB@28_mAd024_2 CB@28_mAd025_1 CB@28_mAd025_2 CB@28_mAd026_1 CB@28_mAd026_2 CB@28_mAd027_1 CB@28_mAd027_2 CB@28_mAd030_1 CB@28_mAd030_2 CB@28_mAd031_1 CB@28_mAd031_2 CB@28_mAd032_1 CB@28_mAd032_2 CB@28_mAd033_1 CB@28_mAd033_2 CB@28_mAd034_1 CB@28_mAd034_2 CB@28_mAd035_1 
+CB@28_mAd035_2 CB@28_mAd036_1 CB@28_mAd036_2 CB@28_mAd037_1 CB@28_mAd037_2 CB@28_mAd040_1 CB@28_mAd040_2 CB@28_mAd041_1 CB@28_mAd041_2 CB@28_mAd042_1 CB@28_mAd042_2 CB@28_mAd043_1 CB@28_mAd043_2 CB@28_mAd044_1 CB@28_mAd044_2 CB@28_mAd045_1 CB@28_mAd045_2 CB@28_mAd046_1 CB@28_mAd046_2 CB@28_mAd047_1 CB@28_mAd047_2 CB@28_mAd050_1 CB@28_mAd050_2 CB@28_mAd051_1 CB@28_mAd051_2 CB@28_mAd052_1 CB@28_mAd052_2 CB@28_mAd053_1 CB@28_mAd053_2 CB@28_mAd054_1 CB@28_mAd054_2 CB@28_mAd055_1 CB@28_mAd055_2 CB@28_mAd056_1 
+CB@28_mAd056_2 CB@28_mAd057_1 CB@28_mAd057_2 CB@28_mAd060_1 CB@28_mAd060_2 CB@28_mAd066_1 CB@28_mAd066_2 CB@28_mAd067_1 CB@28_mAd067_2 CB@28_mAd100_1 CB@28_mAd100_2 CB@28_mAd101_1 CB@28_mAd101_2 CB@28_mAd102_1 CB@28_mAd102_2 CB@28_mAd110_1 CB@28_mAd110_2 CB@28_mAd111_1 CB@28_mAd111_2 CB@28_mAd112_1 CB@28_mAd112_2 CB@28_mAd113_1 CB@28_mAd113_2 CB@28_mAd114_1 CB@28_mAd114_2 CB@28_mAd115_1 CB@28_mAd115_2 CB@28_mAd116_1 CB@28_mAd116_2 CB@28_mAd117_1 CB@28_mAd117_2 CB@28_mAd120_1 CB@28_mAd120_2 CB@28_mAd121_1 
+CB@28_mAd121_2 CB@28_mAd122_1 CB@28_mAd122_2 CB@28_mAd123_1 CB@28_mAd123_2 CB@28_mAd124_1 CB@28_mAd124_2 CB@28_mAd125_1 CB@28_mAd125_2 CB@28_mAd126_1 CB@28_mAd126_2 CB@28_mAd127_1 CB@28_mAd127_2 CB@28_mAd130_1 CB@28_mAd130_2 CB@28_mAd131_1 CB@28_mAd131_2 CB@28_mAd132_1 CB@28_mAd132_2 CB@28_mAd133_1 CB@28_mAd133_2 CB@28_mAd134_1 CB@28_mAd134_2 CB@28_mAd135_1 CB@28_mAd135_2 CB@28_mAd136_1 CB@28_mAd136_2 CB@28_mAd137_1 CB@28_mAd137_2 CB@28_mAd140_1 CB@28_mAd140_2 CB@28_mAd141_1 CB@28_mAd141_2 CB@28_mAd142_1 
+CB@28_mAd142_2 CB@28_mAd143_1 CB@28_mAd143_2 CB@28_mAd144_1 CB@28_mAd144_2 CB@28_mAd145_1 CB@28_mAd145_2 CB@28_mAd146_1 CB@28_mAd146_2 CB@28_mAd147_1 CB@28_mAd147_2 CB@28_mAd150_1 CB@28_mAd150_2 CB@28_mAd151_1 CB@28_mAd151_2 CB@28_mAd152_1 CB@28_mAd152_2 CB@28_mAd153_1 CB@28_mAd153_2 CB@28_mAd154_1 CB@28_mAd154_2 CB@28_mAd155_1 CB@28_mAd155_2 CB@28_mAd156_1 CB@28_mAd156_2 CB@28_mAd157_1 CB@28_mAd157_2 CB@28_mAd160_1 CB@28_mAd160_2 CB@28_mAd161_1 CB@28_mAd161_2 CB@28_mAd162_1 CB@28_mAd162_2 CB@28_mAd163_1 
+CB@28_mAd163_2 CB@28_mAd164_1 CB@28_mAd164_2 CB@28_mAd165_1 CB@28_mAd165_2 CB@28_mAd166_1 CB@28_mAd166_2 CB@28_mAd167_1 CB@28_mAd167_2 CB@28_mAd170_1 CB@28_mAd170_2 CB@28_mAd171_1 CB@28_mAd171_2 CB@28_mAd172_1 CB@28_mAd172_2 CB@28_mAd173_1 CB@28_mAd173_2 CB@28_mAd175_1 CB@28_mAd175_2 CB@28_mAd176_1 CB@28_mAd176_2 CB@28_mAd177_1 CB@28_mAd177_2 CB@28_mAd200_1 CB@28_mAd200_2 CB@28_mAd201_1 CB@28_mAd201_2 CB@28_mAd202_1 CB@28_mAd202_2 CB@28_mAd204_1 CB@28_mAd204_2 CB@28_mAd205_1 CB@28_mAd205_2 CB@28_mAd206_1 
+CB@28_mAd206_2 CB@28_mAd207_1 CB@28_mAd207_2 CB@28_mAd210_1 CB@28_mAd210_2 CB@28_mAd211_1 CB@28_mAd211_2 CB@28_mAd212_1 CB@28_mAd212_2 CB@28_mAd213_1 CB@28_mAd213_2 CB@28_mAd214_1 CB@28_mAd214_2 CB@28_mAd215_1 CB@28_mAd215_2 CB@28_mAd216_1 CB@28_mAd216_2 CB@28_mAd217_1 CB@28_mAd217_2 CB@28_mAd220_1 CB@28_mAd220_2 CB@28_mAd221_1 CB@28_mAd221_2 CB@28_mAd222_1 CB@28_mAd222_2 CB@28_mAd223_1 CB@28_mAd223_2 CB@28_mAd224_1 CB@28_mAd224_2 CB@28_mAd225_1 CB@28_mAd225_2 CB@28_mAd226_1 CB@28_mAd226_2 CB@28_mAd227_1 
+CB@28_mAd227_2 CB@28_mAd230_1 CB@28_mAd230_2 CB@28_mAd231_1 CB@28_mAd231_2 CB@28_mAd232_1 CB@28_mAd232_2 CB@28_mAd233_1 CB@28_mAd233_2 CB@28_mAd234_1 CB@28_mAd234_2 CB@28_mAd235_1 CB@28_mAd235_2 CB@28_mAd236_1 CB@28_mAd236_2 CB@28_mAd237_1 CB@28_mAd237_2 CB@28_mAd240_1 CB@28_mAd240_2 CB@28_mAd241_1 CB@28_mAd241_2 CB@28_mAd242_1 CB@28_mAd242_2 CB@28_mAd243_1 CB@28_mAd243_2 CB@28_mAd244_1 CB@28_mAd244_2 CB@28_mAd245_1 CB@28_mAd245_2 CB@28_mAd246_1 CB@28_mAd246_2 CB@28_mAd247_1 CB@28_mAd247_2 CB@28_mAd250_1 
+CB@28_mAd250_2 CB@28_mAd251_1 CB@28_mAd251_2 CB@28_mAd252_1 CB@28_mAd252_2 CB@28_mAd253_1 CB@28_mAd253_2 CB@28_mAd254_1 CB@28_mAd254_2 CB@28_mAd255_1 CB@28_mAd255_2 CB@28_mAd256_1 CB@28_mAd256_2 CB@28_mAd257_1 CB@28_mAd257_2 CB@28_mAd260_1 CB@28_mAd260_2 CB@28_mAd261_1 CB@28_mAd261_2 CB@28_mAd262_1 CB@28_mAd262_2 CB@28_mAd263_1 CB@28_mAd263_2 CB@28_mAd264_1 CB@28_mAd264_2 CB@28_mAd265_1 CB@28_mAd265_2 CB@28_mAd266_1 CB@28_mAd266_2 CB@28_mAd267_1 CB@28_mAd267_2 CB@28_mAd275_1 CB@28_mAd275_2 CB@28_mAd276_1 
+CB@28_mAd276_2 CB@28_mAd277_1 CB@28_mAd277_2 CB@28_mAd300_1 CB@28_mAd300_2 CB@28_mAd310_1 CB@28_mAd310_2 CB@28_mAd311_1 CB@28_mAd311_2 CB@28_mAd317_1 CB@28_mAd317_2 CB@28_mAd320_1 CB@28_mAd320_2 CB@28_mAd321_1 CB@28_mAd321_2 CB@28_mAd322_1 CB@28_mAd322_2 CB@28_mAd323_1 CB@28_mAd323_2 CB@28_mAd324_1 CB@28_mAd324_2 CB@28_mAd325_1 CB@28_mAd325_2 CB@28_mAd326_1 CB@28_mAd326_2 CB@28_mAd327_1 CB@28_mAd327_2 CB@28_mAd330_1 CB@28_mAd330_2 CB@28_mAd331_1 CB@28_mAd331_2 CB@28_mAd332_1 CB@28_mAd332_2 CB@28_mAd333_1 
+CB@28_mAd333_2 CB@28_mAd334_1 CB@28_mAd334_2 CB@28_mAd335_1 CB@28_mAd335_2 CB@28_mAd336_1 CB@28_mAd336_2 CB@28_mAd337_1 CB@28_mAd337_2 CB@28_mAd340_1 CB@28_mAd340_2 CB@28_mAd341_1 CB@28_mAd341_2 CB@28_mAd342_1 CB@28_mAd342_2 CB@28_mAd343_1 CB@28_mAd343_2 CB@28_mAd344_1 CB@28_mAd344_2 CB@28_mAd345_1 CB@28_mAd345_2 CB@28_mAd346_1 CB@28_mAd346_2 CB@28_mAd347_1 CB@28_mAd347_2 CB@28_mAd350_1 CB@28_mAd350_2 CB@28_mAd351_1 CB@28_mAd351_2 CB@28_mAd352_1 CB@28_mAd352_2 CB@28_mAd353_1 CB@28_mAd353_2 CB@28_mAd354_1 
+CB@28_mAd354_2 CB@28_mAd355_1 CB@28_mAd355_2 CB@28_mAd356_1 CB@28_mAd356_2 CB@28_mAd357_1 CB@28_mAd357_2 CB@28_mAd360_1 CB@28_mAd360_2 CB@28_mAd361_1 CB@28_mAd361_2 CB@28_mAd362_1 CB@28_mAd362_2 CB@28_mAd363_1 CB@28_mAd363_2 CB@28_mAd364_1 CB@28_mAd364_2 CB@28_mAd365_1 CB@28_mAd365_2 CB@28_mAd366_1 CB@28_mAd366_2 CB@28_mAd367_1 CB@28_mAd367_2 CB@28_mAd371_1 CB@28_mAd371_2 CB@28_mAd372_1 CB@28_mAd372_2 CB@28_mAd373_1 CB@28_mAd373_2 CB@28_mAd374_1 CB@28_mAd374_2 CB@28_mAd375_1 CB@28_mAd375_2 CB@28_mAd376_1 
+CB@28_mAd376_2 CB@28_mAd377_1 CB@28_mAd377_2 CB@28_mAd400_1 CB@28_mAd400_2 CB@28_mAd401_1 CB@28_mAd401_2 CB@28_mAd402_1 CB@28_mAd402_2 CB@28_mAd403_1 CB@28_mAd403_2 CB@28_mAd404_1 CB@28_mAd404_2 CB@28_mAd405_1 CB@28_mAd405_2 CB@28_mAd406_1 CB@28_mAd406_2 CB@28_mAd407_1 CB@28_mAd407_2 CB@28_mAd410_1 CB@28_mAd410_2 CB@28_mAd411_1 CB@28_mAd411_2 CB@28_mAd412_1 CB@28_mAd412_2 CB@28_mAd413_1 CB@28_mAd413_2 CB@28_mAd414_1 CB@28_mAd414_2 CB@28_mAd415_1 CB@28_mAd415_2 CB@28_mAd416_1 CB@28_mAd416_2 CB@28_mAd417_1 
+CB@28_mAd417_2 CB@28_mAd420_1 CB@28_mAd420_2 CB@28_mAd421_1 CB@28_mAd421_2 CB@28_mAd422_1 CB@28_mAd422_2 CB@28_mAd423_1 CB@28_mAd423_2 CB@28_mAd424_1 CB@28_mAd424_2 CB@28_mAd425_1 CB@28_mAd425_2 CB@28_mAd426_1 CB@28_mAd426_2 CB@28_mAd427_1 CB@28_mAd427_2 CB@28_mAd430_1 CB@28_mAd430_2 CB@28_mAd431_1 CB@28_mAd431_2 CB@28_mAd432_1 CB@28_mAd432_2 CB@28_mAd433_1 CB@28_mAd433_2 CB@28_mAd434_1 CB@28_mAd434_2 CB@28_mAd435_1 CB@28_mAd435_2 CB@28_mAd436_1 CB@28_mAd436_2 CB@28_mAd437_1 CB@28_mAd437_2 CB@28_mAd440_1 
+CB@28_mAd440_2 CB@28_mAd441_1 CB@28_mAd441_2 CB@28_mAd442_1 CB@28_mAd442_2 CB@28_mAd443_1 CB@28_mAd443_2 CB@28_mAd444_1 CB@28_mAd444_2 CB@28_mAd445_1 CB@28_mAd445_2 CB@28_mAd446_1 CB@28_mAd446_2 CB@28_mAd447_1 CB@28_mAd447_2 CB@28_mAd450_1 CB@28_mAd450_2 CB@28_mAd451_1 CB@28_mAd451_2 CB@28_mAd452_1 CB@28_mAd452_2 CB@28_mAd453_1 CB@28_mAd453_2 CB@28_mAd454_1 CB@28_mAd454_2 CB@28_mAd455_1 CB@28_mAd455_2 CB@28_mAd456_1 CB@28_mAd456_2 CB@28_mAd457_1 CB@28_mAd457_2 CB@28_mAd460_1 CB@28_mAd460_2 CB@28_mAd466_1 
+CB@28_mAd466_2 CB@28_mAd467_1 CB@28_mAd467_2 CB@28_mAd500_1 CB@28_mAd500_2 CB@28_mAd501_1 CB@28_mAd501_2 CB@28_mAd502_1 CB@28_mAd502_2 CB@28_mAd508_1 CB@28_mAd508_2 CB@28_mAd509_1 CB@28_mAd509_2 CB@28_mAd512_1 CB@28_mAd512_2 CB@28_mAd513_1 CB@28_mAd513_2 CB@28_mAd514_1 CB@28_mAd514_2 CB@28_mAd515_1 CB@28_mAd515_2 CB@28_mAd516_1 CB@28_mAd516_2 CB@28_mAd517_1 CB@28_mAd517_2 CB@28_mAd520_1 CB@28_mAd520_2 CB@28_mAd521_1 CB@28_mAd521_2 CB@28_mAd522_1 CB@28_mAd522_2 CB@28_mAd523_1 CB@28_mAd523_2 CB@28_mAd524_1 
+CB@28_mAd524_2 CB@28_mAd525_1 CB@28_mAd525_2 CB@28_mAd526_1 CB@28_mAd526_2 CB@28_mAd527_1 CB@28_mAd527_2 CB@28_mAd530_1 CB@28_mAd530_2 CB@28_mAd531_1 CB@28_mAd531_2 CB@28_mAd532_1 CB@28_mAd532_2 CB@28_mAd533_1 CB@28_mAd533_2 CB@28_mAd534_1 CB@28_mAd534_2 CB@28_mAd535_1 CB@28_mAd535_2 CB@28_mAd536_1 CB@28_mAd536_2 CB@28_mAd537_1 CB@28_mAd537_2 CB@28_mAd540_1 CB@28_mAd540_2 CB@28_mAd541_1 CB@28_mAd541_2 CB@28_mAd542_1 CB@28_mAd542_2 CB@28_mAd543_1 CB@28_mAd543_2 CB@28_mAd544_1 CB@28_mAd544_2 CB@28_mAd545_1 
+CB@28_mAd545_2 CB@28_mAd546_1 CB@28_mAd546_2 CB@28_mAd547_1 CB@28_mAd547_2 CB@28_mAd550_1 CB@28_mAd550_2 CB@28_mAd551_1 CB@28_mAd551_2 CB@28_mAd552_1 CB@28_mAd552_2 CB@28_mAd553_1 CB@28_mAd553_2 CB@28_mAd554_1 CB@28_mAd554_2 CB@28_mAd555_1 CB@28_mAd555_2 CB@28_mAd556_1 CB@28_mAd556_2 CB@28_mAd557_1 CB@28_mAd557_2 CB@28_mAd560_1 CB@28_mAd560_2 CB@28_mAd561_1 CB@28_mAd561_2 CB@28_mAd562_1 CB@28_mAd562_2 CB@28_mAd563_1 CB@28_mAd563_2 CB@28_mAd564_1 CB@28_mAd564_2 CB@28_mAd565_1 CB@28_mAd565_2 CB@28_mAd566_1 
+CB@28_mAd566_2 CB@28_mAd567_1 CB@28_mAd567_2 CB@28_mAd570_1 CB@28_mAd570_2 CB@28_mAd571_1 CB@28_mAd571_2 CB@28_mAd572_1 CB@28_mAd572_2 CB@28_mAd573_1 CB@28_mAd573_2 CB@28_mAd575_1 CB@28_mAd575_2 CB@28_mAd576_1 CB@28_mAd576_2 CB@28_mAd577_1 CB@28_mAd577_2 CB@28_mAd600_1 CB@28_mAd600_2 CB@28_mAd601_1 CB@28_mAd601_2 CB@28_mAd602_1 CB@28_mAd602_2 CB@28_mAd604_1 CB@28_mAd604_2 CB@28_mAd605_1 CB@28_mAd605_2 CB@28_mAd606_1 CB@28_mAd606_2 CB@28_mAd607_1 CB@28_mAd607_2 CB@28_mAd610_1 CB@28_mAd610_2 CB@28_mAd611_1 
+CB@28_mAd611_2 CB@28_mAd612_1 CB@28_mAd612_2 CB@28_mAd613_1 CB@28_mAd613_2 CB@28_mAd614_1 CB@28_mAd614_2 CB@28_mAd615_1 CB@28_mAd615_2 CB@28_mAd616_1 CB@28_mAd616_2 CB@28_mAd617_1 CB@28_mAd617_2 CB@28_mAd620_1 CB@28_mAd620_2 CB@28_mAd621_1 CB@28_mAd621_2 CB@28_mAd622_1 CB@28_mAd622_2 CB@28_mAd623_1 CB@28_mAd623_2 CB@28_mAd624_1 CB@28_mAd624_2 CB@28_mAd625_1 CB@28_mAd625_2 CB@28_mAd626_1 CB@28_mAd626_2 CB@28_mAd627_1 CB@28_mAd627_2 CB@28_mAd630_1 CB@28_mAd630_2 CB@28_mAd631_1 CB@28_mAd631_2 CB@28_mAd632_1 
+CB@28_mAd632_2 CB@28_mAd633_1 CB@28_mAd633_2 CB@28_mAd634_1 CB@28_mAd634_2 CB@28_mAd635_1 CB@28_mAd635_2 CB@28_mAd636_1 CB@28_mAd636_2 CB@28_mAd637_1 CB@28_mAd637_2 CB@28_mAd640_1 CB@28_mAd640_2 CB@28_mAd641_1 CB@28_mAd641_2 CB@28_mAd642_1 CB@28_mAd642_2 CB@28_mAd643_1 CB@28_mAd643_2 CB@28_mAd644_1 CB@28_mAd644_2 CB@28_mAd645_1 CB@28_mAd645_2 CB@28_mAd646_1 CB@28_mAd646_2 CB@28_mAd647_1 CB@28_mAd647_2 CB@28_mAd650_1 CB@28_mAd650_2 CB@28_mAd651_1 CB@28_mAd651_2 CB@28_mAd652_1 CB@28_mAd652_2 CB@28_mAd653_1 
+CB@28_mAd653_2 CB@28_mAd654_1 CB@28_mAd654_2 CB@28_mAd655_1 CB@28_mAd655_2 CB@28_mAd656_1 CB@28_mAd656_2 CB@28_mAd657_1 CB@28_mAd657_2 CB@28_mAd660_1 CB@28_mAd660_2 CB@28_mAd661_1 CB@28_mAd661_2 CB@28_mAd662_1 CB@28_mAd662_2 CB@28_mAd663_1 CB@28_mAd663_2 CB@28_mAd664_1 CB@28_mAd664_2 CB@28_mAd665_1 CB@28_mAd665_2 CB@28_mAd666_1 CB@28_mAd666_2 CB@28_mAd667_1 CB@28_mAd667_2 CB@28_mAd675_1 CB@28_mAd675_2 CB@28_mAd676_1 CB@28_mAd676_2 CB@28_mAd677_1 CB@28_mAd677_2 CB@28_mAd700_1 CB@28_mAd700_2 CB@28_mAd710_1 
+CB@28_mAd710_2 CB@28_mAd711_1 CB@28_mAd711_2 CB@28_mAd717_1 CB@28_mAd717_2 CB@28_mAd720_1 CB@28_mAd720_2 CB@28_mAd721_1 CB@28_mAd721_2 CB@28_mAd722_1 CB@28_mAd722_2 CB@28_mAd723_1 CB@28_mAd723_2 CB@28_mAd724_1 CB@28_mAd724_2 CB@28_mAd725_1 CB@28_mAd725_2 CB@28_mAd726_1 CB@28_mAd726_2 CB@28_mAd727_1 CB@28_mAd727_2 CB@28_mAd730_1 CB@28_mAd730_2 CB@28_mAd731_1 CB@28_mAd731_2 CB@28_mAd732_1 CB@28_mAd732_2 CB@28_mAd733_1 CB@28_mAd733_2 CB@28_mAd734_1 CB@28_mAd734_2 CB@28_mAd735_1 CB@28_mAd735_2 CB@28_mAd736_1 
+CB@28_mAd736_2 CB@28_mAd737_1 CB@28_mAd737_2 CB@28_mAd740_1 CB@28_mAd740_2 CB@28_mAd741_1 CB@28_mAd741_2 CB@28_mAd742_1 CB@28_mAd742_2 CB@28_mAd743_1 CB@28_mAd743_2 CB@28_mAd744_1 CB@28_mAd744_2 CB@28_mAd745_1 CB@28_mAd745_2 CB@28_mAd746_1 CB@28_mAd746_2 CB@28_mAd747_1 CB@28_mAd747_2 CB@28_mAd750_1 CB@28_mAd750_2 CB@28_mAd751_1 CB@28_mAd751_2 CB@28_mAd752_1 CB@28_mAd752_2 CB@28_mAd753_1 CB@28_mAd753_2 CB@28_mAd754_1 CB@28_mAd754_2 CB@28_mAd755_1 CB@28_mAd755_2 CB@28_mAd756_1 CB@28_mAd756_2 CB@28_mAd757_1 
+CB@28_mAd757_2 CB@28_mAd760_1 CB@28_mAd760_2 CB@28_mAd761_1 CB@28_mAd761_2 CB@28_mAd762_1 CB@28_mAd762_2 CB@28_mAd763_1 CB@28_mAd763_2 CB@28_mAd764_1 CB@28_mAd764_2 CB@28_mAd765_1 CB@28_mAd765_2 CB@28_mAd766_1 CB@28_mAd766_2 CB@28_mAd767_1 CB@28_mAd767_2 CB@28_mAd771_1 CB@28_mAd771_2 CB@28_mAd772_1 CB@28_mAd772_2 CB@28_mAd773_1 CB@28_mAd773_2 CB@28_mAd774_1 CB@28_mAd774_2 CB@28_mAd775_1 CB@28_mAd775_2 CB@28_mAd776_1 CB@28_mAd776_2 CB@28_mAd777_1 CB@28_mAd777_2 CB@28_X0 CB@28_X1 CB@28_X10 CB@28_X11 
+CB@28_X12 CB@28_X13 CB@28_X2 CB@28_X3 CB@28_X4 CB@28_X5 CB@28_X6 CB@28_X7 CB@28_X8 CB@28_X9 CB@28_Y1 CB@28_Y10 CB@28_Y11 CB@28_Y12 CB@28_Y2 CB@28_Y3 CB@28_Y4 CB@28_Y5 CB@28_Y6 CB@28_Y7 CB@28_Y8 CB@28_Y9 CB@28_Z1 CB@28_Z10 CB@28_Z11 CB@28_Z12 CB@28_Z2 CB@28_Z3 CB@28_Z4 CB@28_Z5 CB@28_Z6 CB@28_Z7 CB@28_Z8 CB@28_Z9 _5400TP094__CB
XCB@29 CB@29_K0 CB@29_K1 CB@29_K10 CB@29_K11 CB@29_K12 CB@29_K13 CB@29_K2 CB@29_K3 CB@29_K4 CB@29_K5 CB@29_K6 CB@29_K7 CB@29_K8 CB@29_K9 CB@29_mAd000_1 CB@29_mAd000_2 CB@29_mAd001_1 CB@29_mAd001_2 CB@29_mAd002_1 CB@29_mAd002_2 CB@29_mAd003_1 CB@29_mAd003_2 CB@29_mAd004_1 CB@29_mAd004_2 CB@29_mAd005_1 CB@29_mAd005_2 CB@29_mAd006_1 CB@29_mAd006_2 CB@29_mAd007_1 CB@29_mAd007_2 CB@29_mAd010_1 CB@29_mAd010_2 CB@29_mAd011_1 CB@29_mAd011_2 CB@29_mAd012_1 CB@29_mAd012_2 CB@29_mAd013_1 CB@29_mAd013_2 CB@29_mAd014_1 
+CB@29_mAd014_2 CB@29_mAd015_1 CB@29_mAd015_2 CB@29_mAd016_1 CB@29_mAd016_2 CB@29_mAd017_1 CB@29_mAd017_2 CB@29_mAd020_1 CB@29_mAd020_2 CB@29_mAd021_1 CB@29_mAd021_2 CB@29_mAd022_1 CB@29_mAd022_2 CB@29_mAd023_1 CB@29_mAd023_2 CB@29_mAd024_1 CB@29_mAd024_2 CB@29_mAd025_1 CB@29_mAd025_2 CB@29_mAd026_1 CB@29_mAd026_2 CB@29_mAd027_1 CB@29_mAd027_2 CB@29_mAd030_1 CB@29_mAd030_2 CB@29_mAd031_1 CB@29_mAd031_2 CB@29_mAd032_1 CB@29_mAd032_2 CB@29_mAd033_1 CB@29_mAd033_2 CB@29_mAd034_1 CB@29_mAd034_2 CB@29_mAd035_1 
+CB@29_mAd035_2 CB@29_mAd036_1 CB@29_mAd036_2 CB@29_mAd037_1 CB@29_mAd037_2 CB@29_mAd040_1 CB@29_mAd040_2 CB@29_mAd041_1 CB@29_mAd041_2 CB@29_mAd042_1 CB@29_mAd042_2 CB@29_mAd043_1 CB@29_mAd043_2 CB@29_mAd044_1 CB@29_mAd044_2 CB@29_mAd045_1 CB@29_mAd045_2 CB@29_mAd046_1 CB@29_mAd046_2 CB@29_mAd047_1 CB@29_mAd047_2 CB@29_mAd050_1 CB@29_mAd050_2 CB@29_mAd051_1 CB@29_mAd051_2 CB@29_mAd052_1 CB@29_mAd052_2 CB@29_mAd053_1 CB@29_mAd053_2 CB@29_mAd054_1 CB@29_mAd054_2 CB@29_mAd055_1 CB@29_mAd055_2 CB@29_mAd056_1 
+CB@29_mAd056_2 CB@29_mAd057_1 CB@29_mAd057_2 CB@29_mAd060_1 CB@29_mAd060_2 CB@29_mAd066_1 CB@29_mAd066_2 CB@29_mAd067_1 CB@29_mAd067_2 CB@29_mAd100_1 CB@29_mAd100_2 CB@29_mAd101_1 CB@29_mAd101_2 CB@29_mAd102_1 CB@29_mAd102_2 CB@29_mAd110_1 CB@29_mAd110_2 CB@29_mAd111_1 CB@29_mAd111_2 CB@29_mAd112_1 CB@29_mAd112_2 CB@29_mAd113_1 CB@29_mAd113_2 CB@29_mAd114_1 CB@29_mAd114_2 CB@29_mAd115_1 CB@29_mAd115_2 CB@29_mAd116_1 CB@29_mAd116_2 CB@29_mAd117_1 CB@29_mAd117_2 CB@29_mAd120_1 CB@29_mAd120_2 CB@29_mAd121_1 
+CB@29_mAd121_2 CB@29_mAd122_1 CB@29_mAd122_2 CB@29_mAd123_1 CB@29_mAd123_2 CB@29_mAd124_1 CB@29_mAd124_2 CB@29_mAd125_1 CB@29_mAd125_2 CB@29_mAd126_1 CB@29_mAd126_2 CB@29_mAd127_1 CB@29_mAd127_2 CB@29_mAd130_1 CB@29_mAd130_2 CB@29_mAd131_1 CB@29_mAd131_2 CB@29_mAd132_1 CB@29_mAd132_2 CB@29_mAd133_1 CB@29_mAd133_2 CB@29_mAd134_1 CB@29_mAd134_2 CB@29_mAd135_1 CB@29_mAd135_2 CB@29_mAd136_1 CB@29_mAd136_2 CB@29_mAd137_1 CB@29_mAd137_2 CB@29_mAd140_1 CB@29_mAd140_2 CB@29_mAd141_1 CB@29_mAd141_2 CB@29_mAd142_1 
+CB@29_mAd142_2 CB@29_mAd143_1 CB@29_mAd143_2 CB@29_mAd144_1 CB@29_mAd144_2 CB@29_mAd145_1 CB@29_mAd145_2 CB@29_mAd146_1 CB@29_mAd146_2 CB@29_mAd147_1 CB@29_mAd147_2 CB@29_mAd150_1 CB@29_mAd150_2 CB@29_mAd151_1 CB@29_mAd151_2 CB@29_mAd152_1 CB@29_mAd152_2 CB@29_mAd153_1 CB@29_mAd153_2 CB@29_mAd154_1 CB@29_mAd154_2 CB@29_mAd155_1 CB@29_mAd155_2 CB@29_mAd156_1 CB@29_mAd156_2 CB@29_mAd157_1 CB@29_mAd157_2 CB@29_mAd160_1 CB@29_mAd160_2 CB@29_mAd161_1 CB@29_mAd161_2 CB@29_mAd162_1 CB@29_mAd162_2 CB@29_mAd163_1 
+CB@29_mAd163_2 CB@29_mAd164_1 CB@29_mAd164_2 CB@29_mAd165_1 CB@29_mAd165_2 CB@29_mAd166_1 CB@29_mAd166_2 CB@29_mAd167_1 CB@29_mAd167_2 CB@29_mAd170_1 CB@29_mAd170_2 CB@29_mAd171_1 CB@29_mAd171_2 CB@29_mAd172_1 CB@29_mAd172_2 CB@29_mAd173_1 CB@29_mAd173_2 CB@29_mAd175_1 CB@29_mAd175_2 CB@29_mAd176_1 CB@29_mAd176_2 CB@29_mAd177_1 CB@29_mAd177_2 CB@29_mAd200_1 CB@29_mAd200_2 CB@29_mAd201_1 CB@29_mAd201_2 CB@29_mAd202_1 CB@29_mAd202_2 CB@29_mAd204_1 CB@29_mAd204_2 CB@29_mAd205_1 CB@29_mAd205_2 CB@29_mAd206_1 
+CB@29_mAd206_2 CB@29_mAd207_1 CB@29_mAd207_2 CB@29_mAd210_1 CB@29_mAd210_2 CB@29_mAd211_1 CB@29_mAd211_2 CB@29_mAd212_1 CB@29_mAd212_2 CB@29_mAd213_1 CB@29_mAd213_2 CB@29_mAd214_1 CB@29_mAd214_2 CB@29_mAd215_1 CB@29_mAd215_2 CB@29_mAd216_1 CB@29_mAd216_2 CB@29_mAd217_1 CB@29_mAd217_2 CB@29_mAd220_1 CB@29_mAd220_2 CB@29_mAd221_1 CB@29_mAd221_2 CB@29_mAd222_1 CB@29_mAd222_2 CB@29_mAd223_1 CB@29_mAd223_2 CB@29_mAd224_1 CB@29_mAd224_2 CB@29_mAd225_1 CB@29_mAd225_2 CB@29_mAd226_1 CB@29_mAd226_2 CB@29_mAd227_1 
+CB@29_mAd227_2 CB@29_mAd230_1 CB@29_mAd230_2 CB@29_mAd231_1 CB@29_mAd231_2 CB@29_mAd232_1 CB@29_mAd232_2 CB@29_mAd233_1 CB@29_mAd233_2 CB@29_mAd234_1 CB@29_mAd234_2 CB@29_mAd235_1 CB@29_mAd235_2 CB@29_mAd236_1 CB@29_mAd236_2 CB@29_mAd237_1 CB@29_mAd237_2 CB@29_mAd240_1 CB@29_mAd240_2 CB@29_mAd241_1 CB@29_mAd241_2 CB@29_mAd242_1 CB@29_mAd242_2 CB@29_mAd243_1 CB@29_mAd243_2 CB@29_mAd244_1 CB@29_mAd244_2 CB@29_mAd245_1 CB@29_mAd245_2 CB@29_mAd246_1 CB@29_mAd246_2 CB@29_mAd247_1 CB@29_mAd247_2 CB@29_mAd250_1 
+CB@29_mAd250_2 CB@29_mAd251_1 CB@29_mAd251_2 CB@29_mAd252_1 CB@29_mAd252_2 CB@29_mAd253_1 CB@29_mAd253_2 CB@29_mAd254_1 CB@29_mAd254_2 CB@29_mAd255_1 CB@29_mAd255_2 CB@29_mAd256_1 CB@29_mAd256_2 CB@29_mAd257_1 CB@29_mAd257_2 CB@29_mAd260_1 CB@29_mAd260_2 CB@29_mAd261_1 CB@29_mAd261_2 CB@29_mAd262_1 CB@29_mAd262_2 CB@29_mAd263_1 CB@29_mAd263_2 CB@29_mAd264_1 CB@29_mAd264_2 CB@29_mAd265_1 CB@29_mAd265_2 CB@29_mAd266_1 CB@29_mAd266_2 CB@29_mAd267_1 CB@29_mAd267_2 CB@29_mAd275_1 CB@29_mAd275_2 CB@29_mAd276_1 
+CB@29_mAd276_2 CB@29_mAd277_1 CB@29_mAd277_2 CB@29_mAd300_1 CB@29_mAd300_2 CB@29_mAd310_1 CB@29_mAd310_2 CB@29_mAd311_1 CB@29_mAd311_2 CB@29_mAd317_1 CB@29_mAd317_2 CB@29_mAd320_1 CB@29_mAd320_2 CB@29_mAd321_1 CB@29_mAd321_2 CB@29_mAd322_1 CB@29_mAd322_2 CB@29_mAd323_1 CB@29_mAd323_2 CB@29_mAd324_1 CB@29_mAd324_2 CB@29_mAd325_1 CB@29_mAd325_2 CB@29_mAd326_1 CB@29_mAd326_2 CB@29_mAd327_1 CB@29_mAd327_2 CB@29_mAd330_1 CB@29_mAd330_2 CB@29_mAd331_1 CB@29_mAd331_2 CB@29_mAd332_1 CB@29_mAd332_2 CB@29_mAd333_1 
+CB@29_mAd333_2 CB@29_mAd334_1 CB@29_mAd334_2 CB@29_mAd335_1 CB@29_mAd335_2 CB@29_mAd336_1 CB@29_mAd336_2 CB@29_mAd337_1 CB@29_mAd337_2 CB@29_mAd340_1 CB@29_mAd340_2 CB@29_mAd341_1 CB@29_mAd341_2 CB@29_mAd342_1 CB@29_mAd342_2 CB@29_mAd343_1 CB@29_mAd343_2 CB@29_mAd344_1 CB@29_mAd344_2 CB@29_mAd345_1 CB@29_mAd345_2 CB@29_mAd346_1 CB@29_mAd346_2 CB@29_mAd347_1 CB@29_mAd347_2 CB@29_mAd350_1 CB@29_mAd350_2 CB@29_mAd351_1 CB@29_mAd351_2 CB@29_mAd352_1 CB@29_mAd352_2 CB@29_mAd353_1 CB@29_mAd353_2 CB@29_mAd354_1 
+CB@29_mAd354_2 CB@29_mAd355_1 CB@29_mAd355_2 CB@29_mAd356_1 CB@29_mAd356_2 CB@29_mAd357_1 CB@29_mAd357_2 CB@29_mAd360_1 CB@29_mAd360_2 CB@29_mAd361_1 CB@29_mAd361_2 CB@29_mAd362_1 CB@29_mAd362_2 CB@29_mAd363_1 CB@29_mAd363_2 CB@29_mAd364_1 CB@29_mAd364_2 CB@29_mAd365_1 CB@29_mAd365_2 CB@29_mAd366_1 CB@29_mAd366_2 CB@29_mAd367_1 CB@29_mAd367_2 CB@29_mAd371_1 CB@29_mAd371_2 CB@29_mAd372_1 CB@29_mAd372_2 CB@29_mAd373_1 CB@29_mAd373_2 CB@29_mAd374_1 CB@29_mAd374_2 CB@29_mAd375_1 CB@29_mAd375_2 CB@29_mAd376_1 
+CB@29_mAd376_2 CB@29_mAd377_1 CB@29_mAd377_2 CB@29_mAd400_1 CB@29_mAd400_2 CB@29_mAd401_1 CB@29_mAd401_2 CB@29_mAd402_1 CB@29_mAd402_2 CB@29_mAd403_1 CB@29_mAd403_2 CB@29_mAd404_1 CB@29_mAd404_2 CB@29_mAd405_1 CB@29_mAd405_2 CB@29_mAd406_1 CB@29_mAd406_2 CB@29_mAd407_1 CB@29_mAd407_2 CB@29_mAd410_1 CB@29_mAd410_2 CB@29_mAd411_1 CB@29_mAd411_2 CB@29_mAd412_1 CB@29_mAd412_2 CB@29_mAd413_1 CB@29_mAd413_2 CB@29_mAd414_1 CB@29_mAd414_2 CB@29_mAd415_1 CB@29_mAd415_2 CB@29_mAd416_1 CB@29_mAd416_2 CB@29_mAd417_1 
+CB@29_mAd417_2 CB@29_mAd420_1 CB@29_mAd420_2 CB@29_mAd421_1 CB@29_mAd421_2 CB@29_mAd422_1 CB@29_mAd422_2 CB@29_mAd423_1 CB@29_mAd423_2 CB@29_mAd424_1 CB@29_mAd424_2 CB@29_mAd425_1 CB@29_mAd425_2 CB@29_mAd426_1 CB@29_mAd426_2 CB@29_mAd427_1 CB@29_mAd427_2 CB@29_mAd430_1 CB@29_mAd430_2 CB@29_mAd431_1 CB@29_mAd431_2 CB@29_mAd432_1 CB@29_mAd432_2 CB@29_mAd433_1 CB@29_mAd433_2 CB@29_mAd434_1 CB@29_mAd434_2 CB@29_mAd435_1 CB@29_mAd435_2 CB@29_mAd436_1 CB@29_mAd436_2 CB@29_mAd437_1 CB@29_mAd437_2 CB@29_mAd440_1 
+CB@29_mAd440_2 CB@29_mAd441_1 CB@29_mAd441_2 CB@29_mAd442_1 CB@29_mAd442_2 CB@29_mAd443_1 CB@29_mAd443_2 CB@29_mAd444_1 CB@29_mAd444_2 CB@29_mAd445_1 CB@29_mAd445_2 CB@29_mAd446_1 CB@29_mAd446_2 CB@29_mAd447_1 CB@29_mAd447_2 CB@29_mAd450_1 CB@29_mAd450_2 CB@29_mAd451_1 CB@29_mAd451_2 CB@29_mAd452_1 CB@29_mAd452_2 CB@29_mAd453_1 CB@29_mAd453_2 CB@29_mAd454_1 CB@29_mAd454_2 CB@29_mAd455_1 CB@29_mAd455_2 CB@29_mAd456_1 CB@29_mAd456_2 CB@29_mAd457_1 CB@29_mAd457_2 CB@29_mAd460_1 CB@29_mAd460_2 CB@29_mAd466_1 
+CB@29_mAd466_2 CB@29_mAd467_1 CB@29_mAd467_2 CB@29_mAd500_1 CB@29_mAd500_2 CB@29_mAd501_1 CB@29_mAd501_2 CB@29_mAd502_1 CB@29_mAd502_2 CB@29_mAd508_1 CB@29_mAd508_2 CB@29_mAd509_1 CB@29_mAd509_2 CB@29_mAd512_1 CB@29_mAd512_2 CB@29_mAd513_1 CB@29_mAd513_2 CB@29_mAd514_1 CB@29_mAd514_2 CB@29_mAd515_1 CB@29_mAd515_2 CB@29_mAd516_1 CB@29_mAd516_2 CB@29_mAd517_1 CB@29_mAd517_2 CB@29_mAd520_1 CB@29_mAd520_2 CB@29_mAd521_1 CB@29_mAd521_2 CB@29_mAd522_1 CB@29_mAd522_2 CB@29_mAd523_1 CB@29_mAd523_2 CB@29_mAd524_1 
+CB@29_mAd524_2 CB@29_mAd525_1 CB@29_mAd525_2 CB@29_mAd526_1 CB@29_mAd526_2 CB@29_mAd527_1 CB@29_mAd527_2 CB@29_mAd530_1 CB@29_mAd530_2 CB@29_mAd531_1 CB@29_mAd531_2 CB@29_mAd532_1 CB@29_mAd532_2 CB@29_mAd533_1 CB@29_mAd533_2 CB@29_mAd534_1 CB@29_mAd534_2 CB@29_mAd535_1 CB@29_mAd535_2 CB@29_mAd536_1 CB@29_mAd536_2 CB@29_mAd537_1 CB@29_mAd537_2 CB@29_mAd540_1 CB@29_mAd540_2 CB@29_mAd541_1 CB@29_mAd541_2 CB@29_mAd542_1 CB@29_mAd542_2 CB@29_mAd543_1 CB@29_mAd543_2 CB@29_mAd544_1 CB@29_mAd544_2 CB@29_mAd545_1 
+CB@29_mAd545_2 CB@29_mAd546_1 CB@29_mAd546_2 CB@29_mAd547_1 CB@29_mAd547_2 CB@29_mAd550_1 CB@29_mAd550_2 CB@29_mAd551_1 CB@29_mAd551_2 CB@29_mAd552_1 CB@29_mAd552_2 CB@29_mAd553_1 CB@29_mAd553_2 CB@29_mAd554_1 CB@29_mAd554_2 CB@29_mAd555_1 CB@29_mAd555_2 CB@29_mAd556_1 CB@29_mAd556_2 CB@29_mAd557_1 CB@29_mAd557_2 CB@29_mAd560_1 CB@29_mAd560_2 CB@29_mAd561_1 CB@29_mAd561_2 CB@29_mAd562_1 CB@29_mAd562_2 CB@29_mAd563_1 CB@29_mAd563_2 CB@29_mAd564_1 CB@29_mAd564_2 CB@29_mAd565_1 CB@29_mAd565_2 CB@29_mAd566_1 
+CB@29_mAd566_2 CB@29_mAd567_1 CB@29_mAd567_2 CB@29_mAd570_1 CB@29_mAd570_2 CB@29_mAd571_1 CB@29_mAd571_2 CB@29_mAd572_1 CB@29_mAd572_2 CB@29_mAd573_1 CB@29_mAd573_2 CB@29_mAd575_1 CB@29_mAd575_2 CB@29_mAd576_1 CB@29_mAd576_2 CB@29_mAd577_1 CB@29_mAd577_2 CB@29_mAd600_1 CB@29_mAd600_2 CB@29_mAd601_1 CB@29_mAd601_2 CB@29_mAd602_1 CB@29_mAd602_2 CB@29_mAd604_1 CB@29_mAd604_2 CB@29_mAd605_1 CB@29_mAd605_2 CB@29_mAd606_1 CB@29_mAd606_2 CB@29_mAd607_1 CB@29_mAd607_2 CB@29_mAd610_1 CB@29_mAd610_2 CB@29_mAd611_1 
+CB@29_mAd611_2 CB@29_mAd612_1 CB@29_mAd612_2 CB@29_mAd613_1 CB@29_mAd613_2 CB@29_mAd614_1 CB@29_mAd614_2 CB@29_mAd615_1 CB@29_mAd615_2 CB@29_mAd616_1 CB@29_mAd616_2 CB@29_mAd617_1 CB@29_mAd617_2 CB@29_mAd620_1 CB@29_mAd620_2 CB@29_mAd621_1 CB@29_mAd621_2 CB@29_mAd622_1 CB@29_mAd622_2 CB@29_mAd623_1 CB@29_mAd623_2 CB@29_mAd624_1 CB@29_mAd624_2 CB@29_mAd625_1 CB@29_mAd625_2 CB@29_mAd626_1 CB@29_mAd626_2 CB@29_mAd627_1 CB@29_mAd627_2 CB@29_mAd630_1 CB@29_mAd630_2 CB@29_mAd631_1 CB@29_mAd631_2 CB@29_mAd632_1 
+CB@29_mAd632_2 CB@29_mAd633_1 CB@29_mAd633_2 CB@29_mAd634_1 CB@29_mAd634_2 CB@29_mAd635_1 CB@29_mAd635_2 CB@29_mAd636_1 CB@29_mAd636_2 CB@29_mAd637_1 CB@29_mAd637_2 CB@29_mAd640_1 CB@29_mAd640_2 CB@29_mAd641_1 CB@29_mAd641_2 CB@29_mAd642_1 CB@29_mAd642_2 CB@29_mAd643_1 CB@29_mAd643_2 CB@29_mAd644_1 CB@29_mAd644_2 CB@29_mAd645_1 CB@29_mAd645_2 CB@29_mAd646_1 CB@29_mAd646_2 CB@29_mAd647_1 CB@29_mAd647_2 CB@29_mAd650_1 CB@29_mAd650_2 CB@29_mAd651_1 CB@29_mAd651_2 CB@29_mAd652_1 CB@29_mAd652_2 CB@29_mAd653_1 
+CB@29_mAd653_2 CB@29_mAd654_1 CB@29_mAd654_2 CB@29_mAd655_1 CB@29_mAd655_2 CB@29_mAd656_1 CB@29_mAd656_2 CB@29_mAd657_1 CB@29_mAd657_2 CB@29_mAd660_1 CB@29_mAd660_2 CB@29_mAd661_1 CB@29_mAd661_2 CB@29_mAd662_1 CB@29_mAd662_2 CB@29_mAd663_1 CB@29_mAd663_2 CB@29_mAd664_1 CB@29_mAd664_2 CB@29_mAd665_1 CB@29_mAd665_2 CB@29_mAd666_1 CB@29_mAd666_2 CB@29_mAd667_1 CB@29_mAd667_2 CB@29_mAd675_1 CB@29_mAd675_2 CB@29_mAd676_1 CB@29_mAd676_2 CB@29_mAd677_1 CB@29_mAd677_2 CB@29_mAd700_1 CB@29_mAd700_2 CB@29_mAd710_1 
+CB@29_mAd710_2 CB@29_mAd711_1 CB@29_mAd711_2 CB@29_mAd717_1 CB@29_mAd717_2 CB@29_mAd720_1 CB@29_mAd720_2 CB@29_mAd721_1 CB@29_mAd721_2 CB@29_mAd722_1 CB@29_mAd722_2 CB@29_mAd723_1 CB@29_mAd723_2 CB@29_mAd724_1 CB@29_mAd724_2 CB@29_mAd725_1 CB@29_mAd725_2 CB@29_mAd726_1 CB@29_mAd726_2 CB@29_mAd727_1 CB@29_mAd727_2 CB@29_mAd730_1 CB@29_mAd730_2 CB@29_mAd731_1 CB@29_mAd731_2 CB@29_mAd732_1 CB@29_mAd732_2 CB@29_mAd733_1 CB@29_mAd733_2 CB@29_mAd734_1 CB@29_mAd734_2 CB@29_mAd735_1 CB@29_mAd735_2 CB@29_mAd736_1 
+CB@29_mAd736_2 CB@29_mAd737_1 CB@29_mAd737_2 CB@29_mAd740_1 CB@29_mAd740_2 CB@29_mAd741_1 CB@29_mAd741_2 CB@29_mAd742_1 CB@29_mAd742_2 CB@29_mAd743_1 CB@29_mAd743_2 CB@29_mAd744_1 CB@29_mAd744_2 CB@29_mAd745_1 CB@29_mAd745_2 CB@29_mAd746_1 CB@29_mAd746_2 CB@29_mAd747_1 CB@29_mAd747_2 CB@29_mAd750_1 CB@29_mAd750_2 CB@29_mAd751_1 CB@29_mAd751_2 CB@29_mAd752_1 CB@29_mAd752_2 CB@29_mAd753_1 CB@29_mAd753_2 CB@29_mAd754_1 CB@29_mAd754_2 CB@29_mAd755_1 CB@29_mAd755_2 CB@29_mAd756_1 CB@29_mAd756_2 CB@29_mAd757_1 
+CB@29_mAd757_2 CB@29_mAd760_1 CB@29_mAd760_2 CB@29_mAd761_1 CB@29_mAd761_2 CB@29_mAd762_1 CB@29_mAd762_2 CB@29_mAd763_1 CB@29_mAd763_2 CB@29_mAd764_1 CB@29_mAd764_2 CB@29_mAd765_1 CB@29_mAd765_2 CB@29_mAd766_1 CB@29_mAd766_2 CB@29_mAd767_1 CB@29_mAd767_2 CB@29_mAd771_1 CB@29_mAd771_2 CB@29_mAd772_1 CB@29_mAd772_2 CB@29_mAd773_1 CB@29_mAd773_2 CB@29_mAd774_1 CB@29_mAd774_2 CB@29_mAd775_1 CB@29_mAd775_2 CB@29_mAd776_1 CB@29_mAd776_2 CB@29_mAd777_1 CB@29_mAd777_2 CB@29_X0 CB@29_X1 CB@29_X10 CB@29_X11 
+CB@29_X12 CB@29_X13 CB@29_X2 CB@29_X3 CB@29_X4 CB@29_X5 CB@29_X6 CB@29_X7 CB@29_X8 CB@29_X9 CB@29_Y1 CB@29_Y10 CB@29_Y11 CB@29_Y12 CB@29_Y2 CB@29_Y3 CB@29_Y4 CB@29_Y5 CB@29_Y6 CB@29_Y7 CB@29_Y8 CB@29_Y9 CB@29_Z1 CB@29_Z10 CB@29_Z11 CB@29_Z12 CB@29_Z2 CB@29_Z3 CB@29_Z4 CB@29_Z5 CB@29_Z6 CB@29_Z7 CB@29_Z8 CB@29_Z9 _5400TP094__CB
XCB@30 CB@30_K0 CB@30_K1 CB@30_K10 CB@30_K11 CB@30_K12 CB@30_K13 CB@30_K2 CB@30_K3 CB@30_K4 CB@30_K5 CB@30_K6 CB@30_K7 CB@30_K8 CB@30_K9 CB@30_mAd000_1 CB@30_mAd000_2 CB@30_mAd001_1 CB@30_mAd001_2 CB@30_mAd002_1 CB@30_mAd002_2 CB@30_mAd003_1 CB@30_mAd003_2 CB@30_mAd004_1 CB@30_mAd004_2 CB@30_mAd005_1 CB@30_mAd005_2 CB@30_mAd006_1 CB@30_mAd006_2 CB@30_mAd007_1 CB@30_mAd007_2 CB@30_mAd010_1 CB@30_mAd010_2 CB@30_mAd011_1 CB@30_mAd011_2 CB@30_mAd012_1 CB@30_mAd012_2 CB@30_mAd013_1 CB@30_mAd013_2 CB@30_mAd014_1 
+CB@30_mAd014_2 CB@30_mAd015_1 CB@30_mAd015_2 CB@30_mAd016_1 CB@30_mAd016_2 CB@30_mAd017_1 CB@30_mAd017_2 CB@30_mAd020_1 CB@30_mAd020_2 CB@30_mAd021_1 CB@30_mAd021_2 CB@30_mAd022_1 CB@30_mAd022_2 CB@30_mAd023_1 CB@30_mAd023_2 CB@30_mAd024_1 CB@30_mAd024_2 CB@30_mAd025_1 CB@30_mAd025_2 CB@30_mAd026_1 CB@30_mAd026_2 CB@30_mAd027_1 CB@30_mAd027_2 CB@30_mAd030_1 CB@30_mAd030_2 CB@30_mAd031_1 CB@30_mAd031_2 CB@30_mAd032_1 CB@30_mAd032_2 CB@30_mAd033_1 CB@30_mAd033_2 CB@30_mAd034_1 CB@30_mAd034_2 CB@30_mAd035_1 
+CB@30_mAd035_2 CB@30_mAd036_1 CB@30_mAd036_2 CB@30_mAd037_1 CB@30_mAd037_2 CB@30_mAd040_1 CB@30_mAd040_2 CB@30_mAd041_1 CB@30_mAd041_2 CB@30_mAd042_1 CB@30_mAd042_2 CB@30_mAd043_1 CB@30_mAd043_2 CB@30_mAd044_1 CB@30_mAd044_2 CB@30_mAd045_1 CB@30_mAd045_2 CB@30_mAd046_1 CB@30_mAd046_2 CB@30_mAd047_1 CB@30_mAd047_2 CB@30_mAd050_1 CB@30_mAd050_2 CB@30_mAd051_1 CB@30_mAd051_2 CB@30_mAd052_1 CB@30_mAd052_2 CB@30_mAd053_1 CB@30_mAd053_2 CB@30_mAd054_1 CB@30_mAd054_2 CB@30_mAd055_1 CB@30_mAd055_2 CB@30_mAd056_1 
+CB@30_mAd056_2 CB@30_mAd057_1 CB@30_mAd057_2 CB@30_mAd060_1 CB@30_mAd060_2 CB@30_mAd066_1 CB@30_mAd066_2 CB@30_mAd067_1 CB@30_mAd067_2 CB@30_mAd100_1 CB@30_mAd100_2 CB@30_mAd101_1 CB@30_mAd101_2 CB@30_mAd102_1 CB@30_mAd102_2 CB@30_mAd110_1 CB@30_mAd110_2 CB@30_mAd111_1 CB@30_mAd111_2 CB@30_mAd112_1 CB@30_mAd112_2 CB@30_mAd113_1 CB@30_mAd113_2 CB@30_mAd114_1 CB@30_mAd114_2 CB@30_mAd115_1 CB@30_mAd115_2 CB@30_mAd116_1 CB@30_mAd116_2 CB@30_mAd117_1 CB@30_mAd117_2 CB@30_mAd120_1 CB@30_mAd120_2 CB@30_mAd121_1 
+CB@30_mAd121_2 CB@30_mAd122_1 CB@30_mAd122_2 CB@30_mAd123_1 CB@30_mAd123_2 CB@30_mAd124_1 CB@30_mAd124_2 CB@30_mAd125_1 CB@30_mAd125_2 CB@30_mAd126_1 CB@30_mAd126_2 CB@30_mAd127_1 CB@30_mAd127_2 CB@30_mAd130_1 CB@30_mAd130_2 CB@30_mAd131_1 CB@30_mAd131_2 CB@30_mAd132_1 CB@30_mAd132_2 CB@30_mAd133_1 CB@30_mAd133_2 CB@30_mAd134_1 CB@30_mAd134_2 CB@30_mAd135_1 CB@30_mAd135_2 CB@30_mAd136_1 CB@30_mAd136_2 CB@30_mAd137_1 CB@30_mAd137_2 CB@30_mAd140_1 CB@30_mAd140_2 CB@30_mAd141_1 CB@30_mAd141_2 CB@30_mAd142_1 
+CB@30_mAd142_2 CB@30_mAd143_1 CB@30_mAd143_2 CB@30_mAd144_1 CB@30_mAd144_2 CB@30_mAd145_1 CB@30_mAd145_2 CB@30_mAd146_1 CB@30_mAd146_2 CB@30_mAd147_1 CB@30_mAd147_2 CB@30_mAd150_1 CB@30_mAd150_2 CB@30_mAd151_1 CB@30_mAd151_2 CB@30_mAd152_1 CB@30_mAd152_2 CB@30_mAd153_1 CB@30_mAd153_2 CB@30_mAd154_1 CB@30_mAd154_2 CB@30_mAd155_1 CB@30_mAd155_2 CB@30_mAd156_1 CB@30_mAd156_2 CB@30_mAd157_1 CB@30_mAd157_2 CB@30_mAd160_1 CB@30_mAd160_2 CB@30_mAd161_1 CB@30_mAd161_2 CB@30_mAd162_1 CB@30_mAd162_2 CB@30_mAd163_1 
+CB@30_mAd163_2 CB@30_mAd164_1 CB@30_mAd164_2 CB@30_mAd165_1 CB@30_mAd165_2 CB@30_mAd166_1 CB@30_mAd166_2 CB@30_mAd167_1 CB@30_mAd167_2 CB@30_mAd170_1 CB@30_mAd170_2 CB@30_mAd171_1 CB@30_mAd171_2 CB@30_mAd172_1 CB@30_mAd172_2 CB@30_mAd173_1 CB@30_mAd173_2 CB@30_mAd175_1 CB@30_mAd175_2 CB@30_mAd176_1 CB@30_mAd176_2 CB@30_mAd177_1 CB@30_mAd177_2 CB@30_mAd200_1 CB@30_mAd200_2 CB@30_mAd201_1 CB@30_mAd201_2 CB@30_mAd202_1 CB@30_mAd202_2 CB@30_mAd204_1 CB@30_mAd204_2 CB@30_mAd205_1 CB@30_mAd205_2 CB@30_mAd206_1 
+CB@30_mAd206_2 CB@30_mAd207_1 CB@30_mAd207_2 CB@30_mAd210_1 CB@30_mAd210_2 CB@30_mAd211_1 CB@30_mAd211_2 CB@30_mAd212_1 CB@30_mAd212_2 CB@30_mAd213_1 CB@30_mAd213_2 CB@30_mAd214_1 CB@30_mAd214_2 CB@30_mAd215_1 CB@30_mAd215_2 CB@30_mAd216_1 CB@30_mAd216_2 CB@30_mAd217_1 CB@30_mAd217_2 CB@30_mAd220_1 CB@30_mAd220_2 CB@30_mAd221_1 CB@30_mAd221_2 CB@30_mAd222_1 CB@30_mAd222_2 CB@30_mAd223_1 CB@30_mAd223_2 CB@30_mAd224_1 CB@30_mAd224_2 CB@30_mAd225_1 CB@30_mAd225_2 CB@30_mAd226_1 CB@30_mAd226_2 CB@30_mAd227_1 
+CB@30_mAd227_2 CB@30_mAd230_1 CB@30_mAd230_2 CB@30_mAd231_1 CB@30_mAd231_2 CB@30_mAd232_1 CB@30_mAd232_2 CB@30_mAd233_1 CB@30_mAd233_2 CB@30_mAd234_1 CB@30_mAd234_2 CB@30_mAd235_1 CB@30_mAd235_2 CB@30_mAd236_1 CB@30_mAd236_2 CB@30_mAd237_1 CB@30_mAd237_2 CB@30_mAd240_1 CB@30_mAd240_2 CB@30_mAd241_1 CB@30_mAd241_2 CB@30_mAd242_1 CB@30_mAd242_2 CB@30_mAd243_1 CB@30_mAd243_2 CB@30_mAd244_1 CB@30_mAd244_2 CB@30_mAd245_1 CB@30_mAd245_2 CB@30_mAd246_1 CB@30_mAd246_2 CB@30_mAd247_1 CB@30_mAd247_2 CB@30_mAd250_1 
+CB@30_mAd250_2 CB@30_mAd251_1 CB@30_mAd251_2 CB@30_mAd252_1 CB@30_mAd252_2 CB@30_mAd253_1 CB@30_mAd253_2 CB@30_mAd254_1 CB@30_mAd254_2 CB@30_mAd255_1 CB@30_mAd255_2 CB@30_mAd256_1 CB@30_mAd256_2 CB@30_mAd257_1 CB@30_mAd257_2 CB@30_mAd260_1 CB@30_mAd260_2 CB@30_mAd261_1 CB@30_mAd261_2 CB@30_mAd262_1 CB@30_mAd262_2 CB@30_mAd263_1 CB@30_mAd263_2 CB@30_mAd264_1 CB@30_mAd264_2 CB@30_mAd265_1 CB@30_mAd265_2 CB@30_mAd266_1 CB@30_mAd266_2 CB@30_mAd267_1 CB@30_mAd267_2 CB@30_mAd275_1 CB@30_mAd275_2 CB@30_mAd276_1 
+CB@30_mAd276_2 CB@30_mAd277_1 CB@30_mAd277_2 CB@30_mAd300_1 CB@30_mAd300_2 CB@30_mAd310_1 CB@30_mAd310_2 CB@30_mAd311_1 CB@30_mAd311_2 CB@30_mAd317_1 CB@30_mAd317_2 CB@30_mAd320_1 CB@30_mAd320_2 CB@30_mAd321_1 CB@30_mAd321_2 CB@30_mAd322_1 CB@30_mAd322_2 CB@30_mAd323_1 CB@30_mAd323_2 CB@30_mAd324_1 CB@30_mAd324_2 CB@30_mAd325_1 CB@30_mAd325_2 CB@30_mAd326_1 CB@30_mAd326_2 CB@30_mAd327_1 CB@30_mAd327_2 CB@30_mAd330_1 CB@30_mAd330_2 CB@30_mAd331_1 CB@30_mAd331_2 CB@30_mAd332_1 CB@30_mAd332_2 CB@30_mAd333_1 
+CB@30_mAd333_2 CB@30_mAd334_1 CB@30_mAd334_2 CB@30_mAd335_1 CB@30_mAd335_2 CB@30_mAd336_1 CB@30_mAd336_2 CB@30_mAd337_1 CB@30_mAd337_2 CB@30_mAd340_1 CB@30_mAd340_2 CB@30_mAd341_1 CB@30_mAd341_2 CB@30_mAd342_1 CB@30_mAd342_2 CB@30_mAd343_1 CB@30_mAd343_2 CB@30_mAd344_1 CB@30_mAd344_2 CB@30_mAd345_1 CB@30_mAd345_2 CB@30_mAd346_1 CB@30_mAd346_2 CB@30_mAd347_1 CB@30_mAd347_2 CB@30_mAd350_1 CB@30_mAd350_2 CB@30_mAd351_1 CB@30_mAd351_2 CB@30_mAd352_1 CB@30_mAd352_2 CB@30_mAd353_1 CB@30_mAd353_2 CB@30_mAd354_1 
+CB@30_mAd354_2 CB@30_mAd355_1 CB@30_mAd355_2 CB@30_mAd356_1 CB@30_mAd356_2 CB@30_mAd357_1 CB@30_mAd357_2 CB@30_mAd360_1 CB@30_mAd360_2 CB@30_mAd361_1 CB@30_mAd361_2 CB@30_mAd362_1 CB@30_mAd362_2 CB@30_mAd363_1 CB@30_mAd363_2 CB@30_mAd364_1 CB@30_mAd364_2 CB@30_mAd365_1 CB@30_mAd365_2 CB@30_mAd366_1 CB@30_mAd366_2 CB@30_mAd367_1 CB@30_mAd367_2 CB@30_mAd371_1 CB@30_mAd371_2 CB@30_mAd372_1 CB@30_mAd372_2 CB@30_mAd373_1 CB@30_mAd373_2 CB@30_mAd374_1 CB@30_mAd374_2 CB@30_mAd375_1 CB@30_mAd375_2 CB@30_mAd376_1 
+CB@30_mAd376_2 CB@30_mAd377_1 CB@30_mAd377_2 CB@30_mAd400_1 CB@30_mAd400_2 CB@30_mAd401_1 CB@30_mAd401_2 CB@30_mAd402_1 CB@30_mAd402_2 CB@30_mAd403_1 CB@30_mAd403_2 CB@30_mAd404_1 CB@30_mAd404_2 CB@30_mAd405_1 CB@30_mAd405_2 CB@30_mAd406_1 CB@30_mAd406_2 CB@30_mAd407_1 CB@30_mAd407_2 CB@30_mAd410_1 CB@30_mAd410_2 CB@30_mAd411_1 CB@30_mAd411_2 CB@30_mAd412_1 CB@30_mAd412_2 CB@30_mAd413_1 CB@30_mAd413_2 CB@30_mAd414_1 CB@30_mAd414_2 CB@30_mAd415_1 CB@30_mAd415_2 CB@30_mAd416_1 CB@30_mAd416_2 CB@30_mAd417_1 
+CB@30_mAd417_2 CB@30_mAd420_1 CB@30_mAd420_2 CB@30_mAd421_1 CB@30_mAd421_2 CB@30_mAd422_1 CB@30_mAd422_2 CB@30_mAd423_1 CB@30_mAd423_2 CB@30_mAd424_1 CB@30_mAd424_2 CB@30_mAd425_1 CB@30_mAd425_2 CB@30_mAd426_1 CB@30_mAd426_2 CB@30_mAd427_1 CB@30_mAd427_2 CB@30_mAd430_1 CB@30_mAd430_2 CB@30_mAd431_1 CB@30_mAd431_2 CB@30_mAd432_1 CB@30_mAd432_2 CB@30_mAd433_1 CB@30_mAd433_2 CB@30_mAd434_1 CB@30_mAd434_2 CB@30_mAd435_1 CB@30_mAd435_2 CB@30_mAd436_1 CB@30_mAd436_2 CB@30_mAd437_1 CB@30_mAd437_2 CB@30_mAd440_1 
+CB@30_mAd440_2 CB@30_mAd441_1 CB@30_mAd441_2 CB@30_mAd442_1 CB@30_mAd442_2 CB@30_mAd443_1 CB@30_mAd443_2 CB@30_mAd444_1 CB@30_mAd444_2 CB@30_mAd445_1 CB@30_mAd445_2 CB@30_mAd446_1 CB@30_mAd446_2 CB@30_mAd447_1 CB@30_mAd447_2 CB@30_mAd450_1 CB@30_mAd450_2 CB@30_mAd451_1 CB@30_mAd451_2 CB@30_mAd452_1 CB@30_mAd452_2 CB@30_mAd453_1 CB@30_mAd453_2 CB@30_mAd454_1 CB@30_mAd454_2 CB@30_mAd455_1 CB@30_mAd455_2 CB@30_mAd456_1 CB@30_mAd456_2 CB@30_mAd457_1 CB@30_mAd457_2 CB@30_mAd460_1 CB@30_mAd460_2 CB@30_mAd466_1 
+CB@30_mAd466_2 CB@30_mAd467_1 CB@30_mAd467_2 CB@30_mAd500_1 CB@30_mAd500_2 CB@30_mAd501_1 CB@30_mAd501_2 CB@30_mAd502_1 CB@30_mAd502_2 CB@30_mAd508_1 CB@30_mAd508_2 CB@30_mAd509_1 CB@30_mAd509_2 CB@30_mAd512_1 CB@30_mAd512_2 CB@30_mAd513_1 CB@30_mAd513_2 CB@30_mAd514_1 CB@30_mAd514_2 CB@30_mAd515_1 CB@30_mAd515_2 CB@30_mAd516_1 CB@30_mAd516_2 CB@30_mAd517_1 CB@30_mAd517_2 CB@30_mAd520_1 CB@30_mAd520_2 CB@30_mAd521_1 CB@30_mAd521_2 CB@30_mAd522_1 CB@30_mAd522_2 CB@30_mAd523_1 CB@30_mAd523_2 CB@30_mAd524_1 
+CB@30_mAd524_2 CB@30_mAd525_1 CB@30_mAd525_2 CB@30_mAd526_1 CB@30_mAd526_2 CB@30_mAd527_1 CB@30_mAd527_2 CB@30_mAd530_1 CB@30_mAd530_2 CB@30_mAd531_1 CB@30_mAd531_2 CB@30_mAd532_1 CB@30_mAd532_2 CB@30_mAd533_1 CB@30_mAd533_2 CB@30_mAd534_1 CB@30_mAd534_2 CB@30_mAd535_1 CB@30_mAd535_2 CB@30_mAd536_1 CB@30_mAd536_2 CB@30_mAd537_1 CB@30_mAd537_2 CB@30_mAd540_1 CB@30_mAd540_2 CB@30_mAd541_1 CB@30_mAd541_2 CB@30_mAd542_1 CB@30_mAd542_2 CB@30_mAd543_1 CB@30_mAd543_2 CB@30_mAd544_1 CB@30_mAd544_2 CB@30_mAd545_1 
+CB@30_mAd545_2 CB@30_mAd546_1 CB@30_mAd546_2 CB@30_mAd547_1 CB@30_mAd547_2 CB@30_mAd550_1 CB@30_mAd550_2 CB@30_mAd551_1 CB@30_mAd551_2 CB@30_mAd552_1 CB@30_mAd552_2 CB@30_mAd553_1 CB@30_mAd553_2 CB@30_mAd554_1 CB@30_mAd554_2 CB@30_mAd555_1 CB@30_mAd555_2 CB@30_mAd556_1 CB@30_mAd556_2 CB@30_mAd557_1 CB@30_mAd557_2 CB@30_mAd560_1 CB@30_mAd560_2 CB@30_mAd561_1 CB@30_mAd561_2 CB@30_mAd562_1 CB@30_mAd562_2 CB@30_mAd563_1 CB@30_mAd563_2 CB@30_mAd564_1 CB@30_mAd564_2 CB@30_mAd565_1 CB@30_mAd565_2 CB@30_mAd566_1 
+CB@30_mAd566_2 CB@30_mAd567_1 CB@30_mAd567_2 CB@30_mAd570_1 CB@30_mAd570_2 CB@30_mAd571_1 CB@30_mAd571_2 CB@30_mAd572_1 CB@30_mAd572_2 CB@30_mAd573_1 CB@30_mAd573_2 CB@30_mAd575_1 CB@30_mAd575_2 CB@30_mAd576_1 CB@30_mAd576_2 CB@30_mAd577_1 CB@30_mAd577_2 CB@30_mAd600_1 CB@30_mAd600_2 CB@30_mAd601_1 CB@30_mAd601_2 CB@30_mAd602_1 CB@30_mAd602_2 CB@30_mAd604_1 CB@30_mAd604_2 CB@30_mAd605_1 CB@30_mAd605_2 CB@30_mAd606_1 CB@30_mAd606_2 CB@30_mAd607_1 CB@30_mAd607_2 CB@30_mAd610_1 CB@30_mAd610_2 CB@30_mAd611_1 
+CB@30_mAd611_2 CB@30_mAd612_1 CB@30_mAd612_2 CB@30_mAd613_1 CB@30_mAd613_2 CB@30_mAd614_1 CB@30_mAd614_2 CB@30_mAd615_1 CB@30_mAd615_2 CB@30_mAd616_1 CB@30_mAd616_2 CB@30_mAd617_1 CB@30_mAd617_2 CB@30_mAd620_1 CB@30_mAd620_2 CB@30_mAd621_1 CB@30_mAd621_2 CB@30_mAd622_1 CB@30_mAd622_2 CB@30_mAd623_1 CB@30_mAd623_2 CB@30_mAd624_1 CB@30_mAd624_2 CB@30_mAd625_1 CB@30_mAd625_2 CB@30_mAd626_1 CB@30_mAd626_2 CB@30_mAd627_1 CB@30_mAd627_2 CB@30_mAd630_1 CB@30_mAd630_2 CB@30_mAd631_1 CB@30_mAd631_2 CB@30_mAd632_1 
+CB@30_mAd632_2 CB@30_mAd633_1 CB@30_mAd633_2 CB@30_mAd634_1 CB@30_mAd634_2 CB@30_mAd635_1 CB@30_mAd635_2 CB@30_mAd636_1 CB@30_mAd636_2 CB@30_mAd637_1 CB@30_mAd637_2 CB@30_mAd640_1 CB@30_mAd640_2 CB@30_mAd641_1 CB@30_mAd641_2 CB@30_mAd642_1 CB@30_mAd642_2 CB@30_mAd643_1 CB@30_mAd643_2 CB@30_mAd644_1 CB@30_mAd644_2 CB@30_mAd645_1 CB@30_mAd645_2 CB@30_mAd646_1 CB@30_mAd646_2 CB@30_mAd647_1 CB@30_mAd647_2 CB@30_mAd650_1 CB@30_mAd650_2 CB@30_mAd651_1 CB@30_mAd651_2 CB@30_mAd652_1 CB@30_mAd652_2 CB@30_mAd653_1 
+CB@30_mAd653_2 CB@30_mAd654_1 CB@30_mAd654_2 CB@30_mAd655_1 CB@30_mAd655_2 CB@30_mAd656_1 CB@30_mAd656_2 CB@30_mAd657_1 CB@30_mAd657_2 CB@30_mAd660_1 CB@30_mAd660_2 CB@30_mAd661_1 CB@30_mAd661_2 CB@30_mAd662_1 CB@30_mAd662_2 CB@30_mAd663_1 CB@30_mAd663_2 CB@30_mAd664_1 CB@30_mAd664_2 CB@30_mAd665_1 CB@30_mAd665_2 CB@30_mAd666_1 CB@30_mAd666_2 CB@30_mAd667_1 CB@30_mAd667_2 CB@30_mAd675_1 CB@30_mAd675_2 CB@30_mAd676_1 CB@30_mAd676_2 CB@30_mAd677_1 CB@30_mAd677_2 CB@30_mAd700_1 CB@30_mAd700_2 CB@30_mAd710_1 
+CB@30_mAd710_2 CB@30_mAd711_1 CB@30_mAd711_2 CB@30_mAd717_1 CB@30_mAd717_2 CB@30_mAd720_1 CB@30_mAd720_2 CB@30_mAd721_1 CB@30_mAd721_2 CB@30_mAd722_1 CB@30_mAd722_2 CB@30_mAd723_1 CB@30_mAd723_2 CB@30_mAd724_1 CB@30_mAd724_2 CB@30_mAd725_1 CB@30_mAd725_2 CB@30_mAd726_1 CB@30_mAd726_2 CB@30_mAd727_1 CB@30_mAd727_2 CB@30_mAd730_1 CB@30_mAd730_2 CB@30_mAd731_1 CB@30_mAd731_2 CB@30_mAd732_1 CB@30_mAd732_2 CB@30_mAd733_1 CB@30_mAd733_2 CB@30_mAd734_1 CB@30_mAd734_2 CB@30_mAd735_1 CB@30_mAd735_2 CB@30_mAd736_1 
+CB@30_mAd736_2 CB@30_mAd737_1 CB@30_mAd737_2 CB@30_mAd740_1 CB@30_mAd740_2 CB@30_mAd741_1 CB@30_mAd741_2 CB@30_mAd742_1 CB@30_mAd742_2 CB@30_mAd743_1 CB@30_mAd743_2 CB@30_mAd744_1 CB@30_mAd744_2 CB@30_mAd745_1 CB@30_mAd745_2 CB@30_mAd746_1 CB@30_mAd746_2 CB@30_mAd747_1 CB@30_mAd747_2 CB@30_mAd750_1 CB@30_mAd750_2 CB@30_mAd751_1 CB@30_mAd751_2 CB@30_mAd752_1 CB@30_mAd752_2 CB@30_mAd753_1 CB@30_mAd753_2 CB@30_mAd754_1 CB@30_mAd754_2 CB@30_mAd755_1 CB@30_mAd755_2 CB@30_mAd756_1 CB@30_mAd756_2 CB@30_mAd757_1 
+CB@30_mAd757_2 CB@30_mAd760_1 CB@30_mAd760_2 CB@30_mAd761_1 CB@30_mAd761_2 CB@30_mAd762_1 CB@30_mAd762_2 CB@30_mAd763_1 CB@30_mAd763_2 CB@30_mAd764_1 CB@30_mAd764_2 CB@30_mAd765_1 CB@30_mAd765_2 CB@30_mAd766_1 CB@30_mAd766_2 CB@30_mAd767_1 CB@30_mAd767_2 CB@30_mAd771_1 CB@30_mAd771_2 CB@30_mAd772_1 CB@30_mAd772_2 CB@30_mAd773_1 CB@30_mAd773_2 CB@30_mAd774_1 CB@30_mAd774_2 CB@30_mAd775_1 CB@30_mAd775_2 CB@30_mAd776_1 CB@30_mAd776_2 CB@30_mAd777_1 CB@30_mAd777_2 CB@30_X0 CB@30_X1 CB@30_X10 CB@30_X11 
+CB@30_X12 CB@30_X13 CB@30_X2 CB@30_X3 CB@30_X4 CB@30_X5 CB@30_X6 CB@30_X7 CB@30_X8 CB@30_X9 CB@30_Y1 CB@30_Y10 CB@30_Y11 CB@30_Y12 CB@30_Y2 CB@30_Y3 CB@30_Y4 CB@30_Y5 CB@30_Y6 CB@30_Y7 CB@30_Y8 CB@30_Y9 CB@30_Z1 CB@30_Z10 CB@30_Z11 CB@30_Z12 CB@30_Z2 CB@30_Z3 CB@30_Z4 CB@30_Z5 CB@30_Z6 CB@30_Z7 CB@30_Z8 CB@30_Z9 _5400TP094__CB
XCB@31 CB@31_K0 CB@31_K1 CB@31_K10 CB@31_K11 CB@31_K12 CB@31_K13 CB@31_K2 CB@31_K3 CB@31_K4 CB@31_K5 CB@31_K6 CB@31_K7 CB@31_K8 CB@31_K9 CB@31_mAd000_1 CB@31_mAd000_2 CB@31_mAd001_1 CB@31_mAd001_2 CB@31_mAd002_1 CB@31_mAd002_2 CB@31_mAd003_1 CB@31_mAd003_2 CB@31_mAd004_1 CB@31_mAd004_2 CB@31_mAd005_1 CB@31_mAd005_2 CB@31_mAd006_1 CB@31_mAd006_2 CB@31_mAd007_1 CB@31_mAd007_2 CB@31_mAd010_1 CB@31_mAd010_2 CB@31_mAd011_1 CB@31_mAd011_2 CB@31_mAd012_1 CB@31_mAd012_2 CB@31_mAd013_1 CB@31_mAd013_2 CB@31_mAd014_1 
+CB@31_mAd014_2 CB@31_mAd015_1 CB@31_mAd015_2 CB@31_mAd016_1 CB@31_mAd016_2 CB@31_mAd017_1 CB@31_mAd017_2 CB@31_mAd020_1 CB@31_mAd020_2 CB@31_mAd021_1 CB@31_mAd021_2 CB@31_mAd022_1 CB@31_mAd022_2 CB@31_mAd023_1 CB@31_mAd023_2 CB@31_mAd024_1 CB@31_mAd024_2 CB@31_mAd025_1 CB@31_mAd025_2 CB@31_mAd026_1 CB@31_mAd026_2 CB@31_mAd027_1 CB@31_mAd027_2 CB@31_mAd030_1 CB@31_mAd030_2 CB@31_mAd031_1 CB@31_mAd031_2 CB@31_mAd032_1 CB@31_mAd032_2 CB@31_mAd033_1 CB@31_mAd033_2 CB@31_mAd034_1 CB@31_mAd034_2 CB@31_mAd035_1 
+CB@31_mAd035_2 CB@31_mAd036_1 CB@31_mAd036_2 CB@31_mAd037_1 CB@31_mAd037_2 CB@31_mAd040_1 CB@31_mAd040_2 CB@31_mAd041_1 CB@31_mAd041_2 CB@31_mAd042_1 CB@31_mAd042_2 CB@31_mAd043_1 CB@31_mAd043_2 CB@31_mAd044_1 CB@31_mAd044_2 CB@31_mAd045_1 CB@31_mAd045_2 CB@31_mAd046_1 CB@31_mAd046_2 CB@31_mAd047_1 CB@31_mAd047_2 CB@31_mAd050_1 CB@31_mAd050_2 CB@31_mAd051_1 CB@31_mAd051_2 CB@31_mAd052_1 CB@31_mAd052_2 CB@31_mAd053_1 CB@31_mAd053_2 CB@31_mAd054_1 CB@31_mAd054_2 CB@31_mAd055_1 CB@31_mAd055_2 CB@31_mAd056_1 
+CB@31_mAd056_2 CB@31_mAd057_1 CB@31_mAd057_2 CB@31_mAd060_1 CB@31_mAd060_2 CB@31_mAd066_1 CB@31_mAd066_2 CB@31_mAd067_1 CB@31_mAd067_2 CB@31_mAd100_1 CB@31_mAd100_2 CB@31_mAd101_1 CB@31_mAd101_2 CB@31_mAd102_1 CB@31_mAd102_2 CB@31_mAd110_1 CB@31_mAd110_2 CB@31_mAd111_1 CB@31_mAd111_2 CB@31_mAd112_1 CB@31_mAd112_2 CB@31_mAd113_1 CB@31_mAd113_2 CB@31_mAd114_1 CB@31_mAd114_2 CB@31_mAd115_1 CB@31_mAd115_2 CB@31_mAd116_1 CB@31_mAd116_2 CB@31_mAd117_1 CB@31_mAd117_2 CB@31_mAd120_1 CB@31_mAd120_2 CB@31_mAd121_1 
+CB@31_mAd121_2 CB@31_mAd122_1 CB@31_mAd122_2 CB@31_mAd123_1 CB@31_mAd123_2 CB@31_mAd124_1 CB@31_mAd124_2 CB@31_mAd125_1 CB@31_mAd125_2 CB@31_mAd126_1 CB@31_mAd126_2 CB@31_mAd127_1 CB@31_mAd127_2 CB@31_mAd130_1 CB@31_mAd130_2 CB@31_mAd131_1 CB@31_mAd131_2 CB@31_mAd132_1 CB@31_mAd132_2 CB@31_mAd133_1 CB@31_mAd133_2 CB@31_mAd134_1 CB@31_mAd134_2 CB@31_mAd135_1 CB@31_mAd135_2 CB@31_mAd136_1 CB@31_mAd136_2 CB@31_mAd137_1 CB@31_mAd137_2 CB@31_mAd140_1 CB@31_mAd140_2 CB@31_mAd141_1 CB@31_mAd141_2 CB@31_mAd142_1 
+CB@31_mAd142_2 CB@31_mAd143_1 CB@31_mAd143_2 CB@31_mAd144_1 CB@31_mAd144_2 CB@31_mAd145_1 CB@31_mAd145_2 CB@31_mAd146_1 CB@31_mAd146_2 CB@31_mAd147_1 CB@31_mAd147_2 CB@31_mAd150_1 CB@31_mAd150_2 CB@31_mAd151_1 CB@31_mAd151_2 CB@31_mAd152_1 CB@31_mAd152_2 CB@31_mAd153_1 CB@31_mAd153_2 CB@31_mAd154_1 CB@31_mAd154_2 CB@31_mAd155_1 CB@31_mAd155_2 CB@31_mAd156_1 CB@31_mAd156_2 CB@31_mAd157_1 CB@31_mAd157_2 CB@31_mAd160_1 CB@31_mAd160_2 CB@31_mAd161_1 CB@31_mAd161_2 CB@31_mAd162_1 CB@31_mAd162_2 CB@31_mAd163_1 
+CB@31_mAd163_2 CB@31_mAd164_1 CB@31_mAd164_2 CB@31_mAd165_1 CB@31_mAd165_2 CB@31_mAd166_1 CB@31_mAd166_2 CB@31_mAd167_1 CB@31_mAd167_2 CB@31_mAd170_1 CB@31_mAd170_2 CB@31_mAd171_1 CB@31_mAd171_2 CB@31_mAd172_1 CB@31_mAd172_2 CB@31_mAd173_1 CB@31_mAd173_2 CB@31_mAd175_1 CB@31_mAd175_2 CB@31_mAd176_1 CB@31_mAd176_2 CB@31_mAd177_1 CB@31_mAd177_2 CB@31_mAd200_1 CB@31_mAd200_2 CB@31_mAd201_1 CB@31_mAd201_2 CB@31_mAd202_1 CB@31_mAd202_2 CB@31_mAd204_1 CB@31_mAd204_2 CB@31_mAd205_1 CB@31_mAd205_2 CB@31_mAd206_1 
+CB@31_mAd206_2 CB@31_mAd207_1 CB@31_mAd207_2 CB@31_mAd210_1 CB@31_mAd210_2 CB@31_mAd211_1 CB@31_mAd211_2 CB@31_mAd212_1 CB@31_mAd212_2 CB@31_mAd213_1 CB@31_mAd213_2 CB@31_mAd214_1 CB@31_mAd214_2 CB@31_mAd215_1 CB@31_mAd215_2 CB@31_mAd216_1 CB@31_mAd216_2 CB@31_mAd217_1 CB@31_mAd217_2 CB@31_mAd220_1 CB@31_mAd220_2 CB@31_mAd221_1 CB@31_mAd221_2 CB@31_mAd222_1 CB@31_mAd222_2 CB@31_mAd223_1 CB@31_mAd223_2 CB@31_mAd224_1 CB@31_mAd224_2 CB@31_mAd225_1 CB@31_mAd225_2 CB@31_mAd226_1 CB@31_mAd226_2 CB@31_mAd227_1 
+CB@31_mAd227_2 CB@31_mAd230_1 CB@31_mAd230_2 CB@31_mAd231_1 CB@31_mAd231_2 CB@31_mAd232_1 CB@31_mAd232_2 CB@31_mAd233_1 CB@31_mAd233_2 CB@31_mAd234_1 CB@31_mAd234_2 CB@31_mAd235_1 CB@31_mAd235_2 CB@31_mAd236_1 CB@31_mAd236_2 CB@31_mAd237_1 CB@31_mAd237_2 CB@31_mAd240_1 CB@31_mAd240_2 CB@31_mAd241_1 CB@31_mAd241_2 CB@31_mAd242_1 CB@31_mAd242_2 CB@31_mAd243_1 CB@31_mAd243_2 CB@31_mAd244_1 CB@31_mAd244_2 CB@31_mAd245_1 CB@31_mAd245_2 CB@31_mAd246_1 CB@31_mAd246_2 CB@31_mAd247_1 CB@31_mAd247_2 CB@31_mAd250_1 
+CB@31_mAd250_2 CB@31_mAd251_1 CB@31_mAd251_2 CB@31_mAd252_1 CB@31_mAd252_2 CB@31_mAd253_1 CB@31_mAd253_2 CB@31_mAd254_1 CB@31_mAd254_2 CB@31_mAd255_1 CB@31_mAd255_2 CB@31_mAd256_1 CB@31_mAd256_2 CB@31_mAd257_1 CB@31_mAd257_2 CB@31_mAd260_1 CB@31_mAd260_2 CB@31_mAd261_1 CB@31_mAd261_2 CB@31_mAd262_1 CB@31_mAd262_2 CB@31_mAd263_1 CB@31_mAd263_2 CB@31_mAd264_1 CB@31_mAd264_2 CB@31_mAd265_1 CB@31_mAd265_2 CB@31_mAd266_1 CB@31_mAd266_2 CB@31_mAd267_1 CB@31_mAd267_2 CB@31_mAd275_1 CB@31_mAd275_2 CB@31_mAd276_1 
+CB@31_mAd276_2 CB@31_mAd277_1 CB@31_mAd277_2 CB@31_mAd300_1 CB@31_mAd300_2 CB@31_mAd310_1 CB@31_mAd310_2 CB@31_mAd311_1 CB@31_mAd311_2 CB@31_mAd317_1 CB@31_mAd317_2 CB@31_mAd320_1 CB@31_mAd320_2 CB@31_mAd321_1 CB@31_mAd321_2 CB@31_mAd322_1 CB@31_mAd322_2 CB@31_mAd323_1 CB@31_mAd323_2 CB@31_mAd324_1 CB@31_mAd324_2 CB@31_mAd325_1 CB@31_mAd325_2 CB@31_mAd326_1 CB@31_mAd326_2 CB@31_mAd327_1 CB@31_mAd327_2 CB@31_mAd330_1 CB@31_mAd330_2 CB@31_mAd331_1 CB@31_mAd331_2 CB@31_mAd332_1 CB@31_mAd332_2 CB@31_mAd333_1 
+CB@31_mAd333_2 CB@31_mAd334_1 CB@31_mAd334_2 CB@31_mAd335_1 CB@31_mAd335_2 CB@31_mAd336_1 CB@31_mAd336_2 CB@31_mAd337_1 CB@31_mAd337_2 CB@31_mAd340_1 CB@31_mAd340_2 CB@31_mAd341_1 CB@31_mAd341_2 CB@31_mAd342_1 CB@31_mAd342_2 CB@31_mAd343_1 CB@31_mAd343_2 CB@31_mAd344_1 CB@31_mAd344_2 CB@31_mAd345_1 CB@31_mAd345_2 CB@31_mAd346_1 CB@31_mAd346_2 CB@31_mAd347_1 CB@31_mAd347_2 CB@31_mAd350_1 CB@31_mAd350_2 CB@31_mAd351_1 CB@31_mAd351_2 CB@31_mAd352_1 CB@31_mAd352_2 CB@31_mAd353_1 CB@31_mAd353_2 CB@31_mAd354_1 
+CB@31_mAd354_2 CB@31_mAd355_1 CB@31_mAd355_2 CB@31_mAd356_1 CB@31_mAd356_2 CB@31_mAd357_1 CB@31_mAd357_2 CB@31_mAd360_1 CB@31_mAd360_2 CB@31_mAd361_1 CB@31_mAd361_2 CB@31_mAd362_1 CB@31_mAd362_2 CB@31_mAd363_1 CB@31_mAd363_2 CB@31_mAd364_1 CB@31_mAd364_2 CB@31_mAd365_1 CB@31_mAd365_2 CB@31_mAd366_1 CB@31_mAd366_2 CB@31_mAd367_1 CB@31_mAd367_2 CB@31_mAd371_1 CB@31_mAd371_2 CB@31_mAd372_1 CB@31_mAd372_2 CB@31_mAd373_1 CB@31_mAd373_2 CB@31_mAd374_1 CB@31_mAd374_2 CB@31_mAd375_1 CB@31_mAd375_2 CB@31_mAd376_1 
+CB@31_mAd376_2 CB@31_mAd377_1 CB@31_mAd377_2 CB@31_mAd400_1 CB@31_mAd400_2 CB@31_mAd401_1 CB@31_mAd401_2 CB@31_mAd402_1 CB@31_mAd402_2 CB@31_mAd403_1 CB@31_mAd403_2 CB@31_mAd404_1 CB@31_mAd404_2 CB@31_mAd405_1 CB@31_mAd405_2 CB@31_mAd406_1 CB@31_mAd406_2 CB@31_mAd407_1 CB@31_mAd407_2 CB@31_mAd410_1 CB@31_mAd410_2 CB@31_mAd411_1 CB@31_mAd411_2 CB@31_mAd412_1 CB@31_mAd412_2 CB@31_mAd413_1 CB@31_mAd413_2 CB@31_mAd414_1 CB@31_mAd414_2 CB@31_mAd415_1 CB@31_mAd415_2 CB@31_mAd416_1 CB@31_mAd416_2 CB@31_mAd417_1 
+CB@31_mAd417_2 CB@31_mAd420_1 CB@31_mAd420_2 CB@31_mAd421_1 CB@31_mAd421_2 CB@31_mAd422_1 CB@31_mAd422_2 CB@31_mAd423_1 CB@31_mAd423_2 CB@31_mAd424_1 CB@31_mAd424_2 CB@31_mAd425_1 CB@31_mAd425_2 CB@31_mAd426_1 CB@31_mAd426_2 CB@31_mAd427_1 CB@31_mAd427_2 CB@31_mAd430_1 CB@31_mAd430_2 CB@31_mAd431_1 CB@31_mAd431_2 CB@31_mAd432_1 CB@31_mAd432_2 CB@31_mAd433_1 CB@31_mAd433_2 CB@31_mAd434_1 CB@31_mAd434_2 CB@31_mAd435_1 CB@31_mAd435_2 CB@31_mAd436_1 CB@31_mAd436_2 CB@31_mAd437_1 CB@31_mAd437_2 CB@31_mAd440_1 
+CB@31_mAd440_2 CB@31_mAd441_1 CB@31_mAd441_2 CB@31_mAd442_1 CB@31_mAd442_2 CB@31_mAd443_1 CB@31_mAd443_2 CB@31_mAd444_1 CB@31_mAd444_2 CB@31_mAd445_1 CB@31_mAd445_2 CB@31_mAd446_1 CB@31_mAd446_2 CB@31_mAd447_1 CB@31_mAd447_2 CB@31_mAd450_1 CB@31_mAd450_2 CB@31_mAd451_1 CB@31_mAd451_2 CB@31_mAd452_1 CB@31_mAd452_2 CB@31_mAd453_1 CB@31_mAd453_2 CB@31_mAd454_1 CB@31_mAd454_2 CB@31_mAd455_1 CB@31_mAd455_2 CB@31_mAd456_1 CB@31_mAd456_2 CB@31_mAd457_1 CB@31_mAd457_2 CB@31_mAd460_1 CB@31_mAd460_2 CB@31_mAd466_1 
+CB@31_mAd466_2 CB@31_mAd467_1 CB@31_mAd467_2 CB@31_mAd500_1 CB@31_mAd500_2 CB@31_mAd501_1 CB@31_mAd501_2 CB@31_mAd502_1 CB@31_mAd502_2 CB@31_mAd508_1 CB@31_mAd508_2 CB@31_mAd509_1 CB@31_mAd509_2 CB@31_mAd512_1 CB@31_mAd512_2 CB@31_mAd513_1 CB@31_mAd513_2 CB@31_mAd514_1 CB@31_mAd514_2 CB@31_mAd515_1 CB@31_mAd515_2 CB@31_mAd516_1 CB@31_mAd516_2 CB@31_mAd517_1 CB@31_mAd517_2 CB@31_mAd520_1 CB@31_mAd520_2 CB@31_mAd521_1 CB@31_mAd521_2 CB@31_mAd522_1 CB@31_mAd522_2 CB@31_mAd523_1 CB@31_mAd523_2 CB@31_mAd524_1 
+CB@31_mAd524_2 CB@31_mAd525_1 CB@31_mAd525_2 CB@31_mAd526_1 CB@31_mAd526_2 CB@31_mAd527_1 CB@31_mAd527_2 CB@31_mAd530_1 CB@31_mAd530_2 CB@31_mAd531_1 CB@31_mAd531_2 CB@31_mAd532_1 CB@31_mAd532_2 CB@31_mAd533_1 CB@31_mAd533_2 CB@31_mAd534_1 CB@31_mAd534_2 CB@31_mAd535_1 CB@31_mAd535_2 CB@31_mAd536_1 CB@31_mAd536_2 CB@31_mAd537_1 CB@31_mAd537_2 CB@31_mAd540_1 CB@31_mAd540_2 CB@31_mAd541_1 CB@31_mAd541_2 CB@31_mAd542_1 CB@31_mAd542_2 CB@31_mAd543_1 CB@31_mAd543_2 CB@31_mAd544_1 CB@31_mAd544_2 CB@31_mAd545_1 
+CB@31_mAd545_2 CB@31_mAd546_1 CB@31_mAd546_2 CB@31_mAd547_1 CB@31_mAd547_2 CB@31_mAd550_1 CB@31_mAd550_2 CB@31_mAd551_1 CB@31_mAd551_2 CB@31_mAd552_1 CB@31_mAd552_2 CB@31_mAd553_1 CB@31_mAd553_2 CB@31_mAd554_1 CB@31_mAd554_2 CB@31_mAd555_1 CB@31_mAd555_2 CB@31_mAd556_1 CB@31_mAd556_2 CB@31_mAd557_1 CB@31_mAd557_2 CB@31_mAd560_1 CB@31_mAd560_2 CB@31_mAd561_1 CB@31_mAd561_2 CB@31_mAd562_1 CB@31_mAd562_2 CB@31_mAd563_1 CB@31_mAd563_2 CB@31_mAd564_1 CB@31_mAd564_2 CB@31_mAd565_1 CB@31_mAd565_2 CB@31_mAd566_1 
+CB@31_mAd566_2 CB@31_mAd567_1 CB@31_mAd567_2 CB@31_mAd570_1 CB@31_mAd570_2 CB@31_mAd571_1 CB@31_mAd571_2 CB@31_mAd572_1 CB@31_mAd572_2 CB@31_mAd573_1 CB@31_mAd573_2 CB@31_mAd575_1 CB@31_mAd575_2 CB@31_mAd576_1 CB@31_mAd576_2 CB@31_mAd577_1 CB@31_mAd577_2 CB@31_mAd600_1 CB@31_mAd600_2 CB@31_mAd601_1 CB@31_mAd601_2 CB@31_mAd602_1 CB@31_mAd602_2 CB@31_mAd604_1 CB@31_mAd604_2 CB@31_mAd605_1 CB@31_mAd605_2 CB@31_mAd606_1 CB@31_mAd606_2 CB@31_mAd607_1 CB@31_mAd607_2 CB@31_mAd610_1 CB@31_mAd610_2 CB@31_mAd611_1 
+CB@31_mAd611_2 CB@31_mAd612_1 CB@31_mAd612_2 CB@31_mAd613_1 CB@31_mAd613_2 CB@31_mAd614_1 CB@31_mAd614_2 CB@31_mAd615_1 CB@31_mAd615_2 CB@31_mAd616_1 CB@31_mAd616_2 CB@31_mAd617_1 CB@31_mAd617_2 CB@31_mAd620_1 CB@31_mAd620_2 CB@31_mAd621_1 CB@31_mAd621_2 CB@31_mAd622_1 CB@31_mAd622_2 CB@31_mAd623_1 CB@31_mAd623_2 CB@31_mAd624_1 CB@31_mAd624_2 CB@31_mAd625_1 CB@31_mAd625_2 CB@31_mAd626_1 CB@31_mAd626_2 CB@31_mAd627_1 CB@31_mAd627_2 CB@31_mAd630_1 CB@31_mAd630_2 CB@31_mAd631_1 CB@31_mAd631_2 CB@31_mAd632_1 
+CB@31_mAd632_2 CB@31_mAd633_1 CB@31_mAd633_2 CB@31_mAd634_1 CB@31_mAd634_2 CB@31_mAd635_1 CB@31_mAd635_2 CB@31_mAd636_1 CB@31_mAd636_2 CB@31_mAd637_1 CB@31_mAd637_2 CB@31_mAd640_1 CB@31_mAd640_2 CB@31_mAd641_1 CB@31_mAd641_2 CB@31_mAd642_1 CB@31_mAd642_2 CB@31_mAd643_1 CB@31_mAd643_2 CB@31_mAd644_1 CB@31_mAd644_2 CB@31_mAd645_1 CB@31_mAd645_2 CB@31_mAd646_1 CB@31_mAd646_2 CB@31_mAd647_1 CB@31_mAd647_2 CB@31_mAd650_1 CB@31_mAd650_2 CB@31_mAd651_1 CB@31_mAd651_2 CB@31_mAd652_1 CB@31_mAd652_2 CB@31_mAd653_1 
+CB@31_mAd653_2 CB@31_mAd654_1 CB@31_mAd654_2 CB@31_mAd655_1 CB@31_mAd655_2 CB@31_mAd656_1 CB@31_mAd656_2 CB@31_mAd657_1 CB@31_mAd657_2 CB@31_mAd660_1 CB@31_mAd660_2 CB@31_mAd661_1 CB@31_mAd661_2 CB@31_mAd662_1 CB@31_mAd662_2 CB@31_mAd663_1 CB@31_mAd663_2 CB@31_mAd664_1 CB@31_mAd664_2 CB@31_mAd665_1 CB@31_mAd665_2 CB@31_mAd666_1 CB@31_mAd666_2 CB@31_mAd667_1 CB@31_mAd667_2 CB@31_mAd675_1 CB@31_mAd675_2 CB@31_mAd676_1 CB@31_mAd676_2 CB@31_mAd677_1 CB@31_mAd677_2 CB@31_mAd700_1 CB@31_mAd700_2 CB@31_mAd710_1 
+CB@31_mAd710_2 CB@31_mAd711_1 CB@31_mAd711_2 CB@31_mAd717_1 CB@31_mAd717_2 CB@31_mAd720_1 CB@31_mAd720_2 CB@31_mAd721_1 CB@31_mAd721_2 CB@31_mAd722_1 CB@31_mAd722_2 CB@31_mAd723_1 CB@31_mAd723_2 CB@31_mAd724_1 CB@31_mAd724_2 CB@31_mAd725_1 CB@31_mAd725_2 CB@31_mAd726_1 CB@31_mAd726_2 CB@31_mAd727_1 CB@31_mAd727_2 CB@31_mAd730_1 CB@31_mAd730_2 CB@31_mAd731_1 CB@31_mAd731_2 CB@31_mAd732_1 CB@31_mAd732_2 CB@31_mAd733_1 CB@31_mAd733_2 CB@31_mAd734_1 CB@31_mAd734_2 CB@31_mAd735_1 CB@31_mAd735_2 CB@31_mAd736_1 
+CB@31_mAd736_2 CB@31_mAd737_1 CB@31_mAd737_2 CB@31_mAd740_1 CB@31_mAd740_2 CB@31_mAd741_1 CB@31_mAd741_2 CB@31_mAd742_1 CB@31_mAd742_2 CB@31_mAd743_1 CB@31_mAd743_2 CB@31_mAd744_1 CB@31_mAd744_2 CB@31_mAd745_1 CB@31_mAd745_2 CB@31_mAd746_1 CB@31_mAd746_2 CB@31_mAd747_1 CB@31_mAd747_2 CB@31_mAd750_1 CB@31_mAd750_2 CB@31_mAd751_1 CB@31_mAd751_2 CB@31_mAd752_1 CB@31_mAd752_2 CB@31_mAd753_1 CB@31_mAd753_2 CB@31_mAd754_1 CB@31_mAd754_2 CB@31_mAd755_1 CB@31_mAd755_2 CB@31_mAd756_1 CB@31_mAd756_2 CB@31_mAd757_1 
+CB@31_mAd757_2 CB@31_mAd760_1 CB@31_mAd760_2 CB@31_mAd761_1 CB@31_mAd761_2 CB@31_mAd762_1 CB@31_mAd762_2 CB@31_mAd763_1 CB@31_mAd763_2 CB@31_mAd764_1 CB@31_mAd764_2 CB@31_mAd765_1 CB@31_mAd765_2 CB@31_mAd766_1 CB@31_mAd766_2 CB@31_mAd767_1 CB@31_mAd767_2 CB@31_mAd771_1 CB@31_mAd771_2 CB@31_mAd772_1 CB@31_mAd772_2 CB@31_mAd773_1 CB@31_mAd773_2 CB@31_mAd774_1 CB@31_mAd774_2 CB@31_mAd775_1 CB@31_mAd775_2 CB@31_mAd776_1 CB@31_mAd776_2 CB@31_mAd777_1 CB@31_mAd777_2 CB@31_X0 CB@31_X1 CB@31_X10 CB@31_X11 
+CB@31_X12 CB@31_X13 CB@31_X2 CB@31_X3 CB@31_X4 CB@31_X5 CB@31_X6 CB@31_X7 CB@31_X8 CB@31_X9 CB@31_Y1 CB@31_Y10 CB@31_Y11 CB@31_Y12 CB@31_Y2 CB@31_Y3 CB@31_Y4 CB@31_Y5 CB@31_Y6 CB@31_Y7 CB@31_Y8 CB@31_Y9 CB@31_Z1 CB@31_Z10 CB@31_Z11 CB@31_Z12 CB@31_Z2 CB@31_Z3 CB@31_Z4 CB@31_Z5 CB@31_Z6 CB@31_Z7 CB@31_Z8 CB@31_Z9 _5400TP094__CB
XCB@32 CB@32_K0 CB@32_K1 CB@32_K10 CB@32_K11 CB@32_K12 CB@32_K13 CB@32_K2 CB@32_K3 CB@32_K4 CB@32_K5 CB@32_K6 CB@32_K7 CB@32_K8 CB@32_K9 CB@32_mAd000_1 CB@32_mAd000_2 CB@32_mAd001_1 CB@32_mAd001_2 CB@32_mAd002_1 CB@32_mAd002_2 CB@32_mAd003_1 CB@32_mAd003_2 CB@32_mAd004_1 CB@32_mAd004_2 CB@32_mAd005_1 CB@32_mAd005_2 CB@32_mAd006_1 CB@32_mAd006_2 CB@32_mAd007_1 CB@32_mAd007_2 CB@32_mAd010_1 CB@32_mAd010_2 CB@32_mAd011_1 CB@32_mAd011_2 CB@32_mAd012_1 CB@32_mAd012_2 CB@32_mAd013_1 CB@32_mAd013_2 CB@32_mAd014_1 
+CB@32_mAd014_2 CB@32_mAd015_1 CB@32_mAd015_2 CB@32_mAd016_1 CB@32_mAd016_2 CB@32_mAd017_1 CB@32_mAd017_2 CB@32_mAd020_1 CB@32_mAd020_2 CB@32_mAd021_1 CB@32_mAd021_2 CB@32_mAd022_1 CB@32_mAd022_2 CB@32_mAd023_1 CB@32_mAd023_2 CB@32_mAd024_1 CB@32_mAd024_2 CB@32_mAd025_1 CB@32_mAd025_2 CB@32_mAd026_1 CB@32_mAd026_2 CB@32_mAd027_1 CB@32_mAd027_2 CB@32_mAd030_1 CB@32_mAd030_2 CB@32_mAd031_1 CB@32_mAd031_2 CB@32_mAd032_1 CB@32_mAd032_2 CB@32_mAd033_1 CB@32_mAd033_2 CB@32_mAd034_1 CB@32_mAd034_2 CB@32_mAd035_1 
+CB@32_mAd035_2 CB@32_mAd036_1 CB@32_mAd036_2 CB@32_mAd037_1 CB@32_mAd037_2 CB@32_mAd040_1 CB@32_mAd040_2 CB@32_mAd041_1 CB@32_mAd041_2 CB@32_mAd042_1 CB@32_mAd042_2 CB@32_mAd043_1 CB@32_mAd043_2 CB@32_mAd044_1 CB@32_mAd044_2 CB@32_mAd045_1 CB@32_mAd045_2 CB@32_mAd046_1 CB@32_mAd046_2 CB@32_mAd047_1 CB@32_mAd047_2 CB@32_mAd050_1 CB@32_mAd050_2 CB@32_mAd051_1 CB@32_mAd051_2 CB@32_mAd052_1 CB@32_mAd052_2 CB@32_mAd053_1 CB@32_mAd053_2 CB@32_mAd054_1 CB@32_mAd054_2 CB@32_mAd055_1 CB@32_mAd055_2 CB@32_mAd056_1 
+CB@32_mAd056_2 CB@32_mAd057_1 CB@32_mAd057_2 CB@32_mAd060_1 CB@32_mAd060_2 CB@32_mAd066_1 CB@32_mAd066_2 CB@32_mAd067_1 CB@32_mAd067_2 CB@32_mAd100_1 CB@32_mAd100_2 CB@32_mAd101_1 CB@32_mAd101_2 CB@32_mAd102_1 CB@32_mAd102_2 CB@32_mAd110_1 CB@32_mAd110_2 CB@32_mAd111_1 CB@32_mAd111_2 CB@32_mAd112_1 CB@32_mAd112_2 CB@32_mAd113_1 CB@32_mAd113_2 CB@32_mAd114_1 CB@32_mAd114_2 CB@32_mAd115_1 CB@32_mAd115_2 CB@32_mAd116_1 CB@32_mAd116_2 CB@32_mAd117_1 CB@32_mAd117_2 CB@32_mAd120_1 CB@32_mAd120_2 CB@32_mAd121_1 
+CB@32_mAd121_2 CB@32_mAd122_1 CB@32_mAd122_2 CB@32_mAd123_1 CB@32_mAd123_2 CB@32_mAd124_1 CB@32_mAd124_2 CB@32_mAd125_1 CB@32_mAd125_2 CB@32_mAd126_1 CB@32_mAd126_2 CB@32_mAd127_1 CB@32_mAd127_2 CB@32_mAd130_1 CB@32_mAd130_2 CB@32_mAd131_1 CB@32_mAd131_2 CB@32_mAd132_1 CB@32_mAd132_2 CB@32_mAd133_1 CB@32_mAd133_2 CB@32_mAd134_1 CB@32_mAd134_2 CB@32_mAd135_1 CB@32_mAd135_2 CB@32_mAd136_1 CB@32_mAd136_2 CB@32_mAd137_1 CB@32_mAd137_2 CB@32_mAd140_1 CB@32_mAd140_2 CB@32_mAd141_1 CB@32_mAd141_2 CB@32_mAd142_1 
+CB@32_mAd142_2 CB@32_mAd143_1 CB@32_mAd143_2 CB@32_mAd144_1 CB@32_mAd144_2 CB@32_mAd145_1 CB@32_mAd145_2 CB@32_mAd146_1 CB@32_mAd146_2 CB@32_mAd147_1 CB@32_mAd147_2 CB@32_mAd150_1 CB@32_mAd150_2 CB@32_mAd151_1 CB@32_mAd151_2 CB@32_mAd152_1 CB@32_mAd152_2 CB@32_mAd153_1 CB@32_mAd153_2 CB@32_mAd154_1 CB@32_mAd154_2 CB@32_mAd155_1 CB@32_mAd155_2 CB@32_mAd156_1 CB@32_mAd156_2 CB@32_mAd157_1 CB@32_mAd157_2 CB@32_mAd160_1 CB@32_mAd160_2 CB@32_mAd161_1 CB@32_mAd161_2 CB@32_mAd162_1 CB@32_mAd162_2 CB@32_mAd163_1 
+CB@32_mAd163_2 CB@32_mAd164_1 CB@32_mAd164_2 CB@32_mAd165_1 CB@32_mAd165_2 CB@32_mAd166_1 CB@32_mAd166_2 CB@32_mAd167_1 CB@32_mAd167_2 CB@32_mAd170_1 CB@32_mAd170_2 CB@32_mAd171_1 CB@32_mAd171_2 CB@32_mAd172_1 CB@32_mAd172_2 CB@32_mAd173_1 CB@32_mAd173_2 CB@32_mAd175_1 CB@32_mAd175_2 CB@32_mAd176_1 CB@32_mAd176_2 CB@32_mAd177_1 CB@32_mAd177_2 CB@32_mAd200_1 CB@32_mAd200_2 CB@32_mAd201_1 CB@32_mAd201_2 CB@32_mAd202_1 CB@32_mAd202_2 CB@32_mAd204_1 CB@32_mAd204_2 CB@32_mAd205_1 CB@32_mAd205_2 CB@32_mAd206_1 
+CB@32_mAd206_2 CB@32_mAd207_1 CB@32_mAd207_2 CB@32_mAd210_1 CB@32_mAd210_2 CB@32_mAd211_1 CB@32_mAd211_2 CB@32_mAd212_1 CB@32_mAd212_2 CB@32_mAd213_1 CB@32_mAd213_2 CB@32_mAd214_1 CB@32_mAd214_2 CB@32_mAd215_1 CB@32_mAd215_2 CB@32_mAd216_1 CB@32_mAd216_2 CB@32_mAd217_1 CB@32_mAd217_2 CB@32_mAd220_1 CB@32_mAd220_2 CB@32_mAd221_1 CB@32_mAd221_2 CB@32_mAd222_1 CB@32_mAd222_2 CB@32_mAd223_1 CB@32_mAd223_2 CB@32_mAd224_1 CB@32_mAd224_2 CB@32_mAd225_1 CB@32_mAd225_2 CB@32_mAd226_1 CB@32_mAd226_2 CB@32_mAd227_1 
+CB@32_mAd227_2 CB@32_mAd230_1 CB@32_mAd230_2 CB@32_mAd231_1 CB@32_mAd231_2 CB@32_mAd232_1 CB@32_mAd232_2 CB@32_mAd233_1 CB@32_mAd233_2 CB@32_mAd234_1 CB@32_mAd234_2 CB@32_mAd235_1 CB@32_mAd235_2 CB@32_mAd236_1 CB@32_mAd236_2 CB@32_mAd237_1 CB@32_mAd237_2 CB@32_mAd240_1 CB@32_mAd240_2 CB@32_mAd241_1 CB@32_mAd241_2 CB@32_mAd242_1 CB@32_mAd242_2 CB@32_mAd243_1 CB@32_mAd243_2 CB@32_mAd244_1 CB@32_mAd244_2 CB@32_mAd245_1 CB@32_mAd245_2 CB@32_mAd246_1 CB@32_mAd246_2 CB@32_mAd247_1 CB@32_mAd247_2 CB@32_mAd250_1 
+CB@32_mAd250_2 CB@32_mAd251_1 CB@32_mAd251_2 CB@32_mAd252_1 CB@32_mAd252_2 CB@32_mAd253_1 CB@32_mAd253_2 CB@32_mAd254_1 CB@32_mAd254_2 CB@32_mAd255_1 CB@32_mAd255_2 CB@32_mAd256_1 CB@32_mAd256_2 CB@32_mAd257_1 CB@32_mAd257_2 CB@32_mAd260_1 CB@32_mAd260_2 CB@32_mAd261_1 CB@32_mAd261_2 CB@32_mAd262_1 CB@32_mAd262_2 CB@32_mAd263_1 CB@32_mAd263_2 CB@32_mAd264_1 CB@32_mAd264_2 CB@32_mAd265_1 CB@32_mAd265_2 CB@32_mAd266_1 CB@32_mAd266_2 CB@32_mAd267_1 CB@32_mAd267_2 CB@32_mAd275_1 CB@32_mAd275_2 CB@32_mAd276_1 
+CB@32_mAd276_2 CB@32_mAd277_1 CB@32_mAd277_2 CB@32_mAd300_1 CB@32_mAd300_2 CB@32_mAd310_1 CB@32_mAd310_2 CB@32_mAd311_1 CB@32_mAd311_2 CB@32_mAd317_1 CB@32_mAd317_2 CB@32_mAd320_1 CB@32_mAd320_2 CB@32_mAd321_1 CB@32_mAd321_2 CB@32_mAd322_1 CB@32_mAd322_2 CB@32_mAd323_1 CB@32_mAd323_2 CB@32_mAd324_1 CB@32_mAd324_2 CB@32_mAd325_1 CB@32_mAd325_2 CB@32_mAd326_1 CB@32_mAd326_2 CB@32_mAd327_1 CB@32_mAd327_2 CB@32_mAd330_1 CB@32_mAd330_2 CB@32_mAd331_1 CB@32_mAd331_2 CB@32_mAd332_1 CB@32_mAd332_2 CB@32_mAd333_1 
+CB@32_mAd333_2 CB@32_mAd334_1 CB@32_mAd334_2 CB@32_mAd335_1 CB@32_mAd335_2 CB@32_mAd336_1 CB@32_mAd336_2 CB@32_mAd337_1 CB@32_mAd337_2 CB@32_mAd340_1 CB@32_mAd340_2 CB@32_mAd341_1 CB@32_mAd341_2 CB@32_mAd342_1 CB@32_mAd342_2 CB@32_mAd343_1 CB@32_mAd343_2 CB@32_mAd344_1 CB@32_mAd344_2 CB@32_mAd345_1 CB@32_mAd345_2 CB@32_mAd346_1 CB@32_mAd346_2 CB@32_mAd347_1 CB@32_mAd347_2 CB@32_mAd350_1 CB@32_mAd350_2 CB@32_mAd351_1 CB@32_mAd351_2 CB@32_mAd352_1 CB@32_mAd352_2 CB@32_mAd353_1 CB@32_mAd353_2 CB@32_mAd354_1 
+CB@32_mAd354_2 CB@32_mAd355_1 CB@32_mAd355_2 CB@32_mAd356_1 CB@32_mAd356_2 CB@32_mAd357_1 CB@32_mAd357_2 CB@32_mAd360_1 CB@32_mAd360_2 CB@32_mAd361_1 CB@32_mAd361_2 CB@32_mAd362_1 CB@32_mAd362_2 CB@32_mAd363_1 CB@32_mAd363_2 CB@32_mAd364_1 CB@32_mAd364_2 CB@32_mAd365_1 CB@32_mAd365_2 CB@32_mAd366_1 CB@32_mAd366_2 CB@32_mAd367_1 CB@32_mAd367_2 CB@32_mAd371_1 CB@32_mAd371_2 CB@32_mAd372_1 CB@32_mAd372_2 CB@32_mAd373_1 CB@32_mAd373_2 CB@32_mAd374_1 CB@32_mAd374_2 CB@32_mAd375_1 CB@32_mAd375_2 CB@32_mAd376_1 
+CB@32_mAd376_2 CB@32_mAd377_1 CB@32_mAd377_2 CB@32_mAd400_1 CB@32_mAd400_2 CB@32_mAd401_1 CB@32_mAd401_2 CB@32_mAd402_1 CB@32_mAd402_2 CB@32_mAd403_1 CB@32_mAd403_2 CB@32_mAd404_1 CB@32_mAd404_2 CB@32_mAd405_1 CB@32_mAd405_2 CB@32_mAd406_1 CB@32_mAd406_2 CB@32_mAd407_1 CB@32_mAd407_2 CB@32_mAd410_1 CB@32_mAd410_2 CB@32_mAd411_1 CB@32_mAd411_2 CB@32_mAd412_1 CB@32_mAd412_2 CB@32_mAd413_1 CB@32_mAd413_2 CB@32_mAd414_1 CB@32_mAd414_2 CB@32_mAd415_1 CB@32_mAd415_2 CB@32_mAd416_1 CB@32_mAd416_2 CB@32_mAd417_1 
+CB@32_mAd417_2 CB@32_mAd420_1 CB@32_mAd420_2 CB@32_mAd421_1 CB@32_mAd421_2 CB@32_mAd422_1 CB@32_mAd422_2 CB@32_mAd423_1 CB@32_mAd423_2 CB@32_mAd424_1 CB@32_mAd424_2 CB@32_mAd425_1 CB@32_mAd425_2 CB@32_mAd426_1 CB@32_mAd426_2 CB@32_mAd427_1 CB@32_mAd427_2 CB@32_mAd430_1 CB@32_mAd430_2 CB@32_mAd431_1 CB@32_mAd431_2 CB@32_mAd432_1 CB@32_mAd432_2 CB@32_mAd433_1 CB@32_mAd433_2 CB@32_mAd434_1 CB@32_mAd434_2 CB@32_mAd435_1 CB@32_mAd435_2 CB@32_mAd436_1 CB@32_mAd436_2 CB@32_mAd437_1 CB@32_mAd437_2 CB@32_mAd440_1 
+CB@32_mAd440_2 CB@32_mAd441_1 CB@32_mAd441_2 CB@32_mAd442_1 CB@32_mAd442_2 CB@32_mAd443_1 CB@32_mAd443_2 CB@32_mAd444_1 CB@32_mAd444_2 CB@32_mAd445_1 CB@32_mAd445_2 CB@32_mAd446_1 CB@32_mAd446_2 CB@32_mAd447_1 CB@32_mAd447_2 CB@32_mAd450_1 CB@32_mAd450_2 CB@32_mAd451_1 CB@32_mAd451_2 CB@32_mAd452_1 CB@32_mAd452_2 CB@32_mAd453_1 CB@32_mAd453_2 CB@32_mAd454_1 CB@32_mAd454_2 CB@32_mAd455_1 CB@32_mAd455_2 CB@32_mAd456_1 CB@32_mAd456_2 CB@32_mAd457_1 CB@32_mAd457_2 CB@32_mAd460_1 CB@32_mAd460_2 CB@32_mAd466_1 
+CB@32_mAd466_2 CB@32_mAd467_1 CB@32_mAd467_2 CB@32_mAd500_1 CB@32_mAd500_2 CB@32_mAd501_1 CB@32_mAd501_2 CB@32_mAd502_1 CB@32_mAd502_2 CB@32_mAd508_1 CB@32_mAd508_2 CB@32_mAd509_1 CB@32_mAd509_2 CB@32_mAd512_1 CB@32_mAd512_2 CB@32_mAd513_1 CB@32_mAd513_2 CB@32_mAd514_1 CB@32_mAd514_2 CB@32_mAd515_1 CB@32_mAd515_2 CB@32_mAd516_1 CB@32_mAd516_2 CB@32_mAd517_1 CB@32_mAd517_2 CB@32_mAd520_1 CB@32_mAd520_2 CB@32_mAd521_1 CB@32_mAd521_2 CB@32_mAd522_1 CB@32_mAd522_2 CB@32_mAd523_1 CB@32_mAd523_2 CB@32_mAd524_1 
+CB@32_mAd524_2 CB@32_mAd525_1 CB@32_mAd525_2 CB@32_mAd526_1 CB@32_mAd526_2 CB@32_mAd527_1 CB@32_mAd527_2 CB@32_mAd530_1 CB@32_mAd530_2 CB@32_mAd531_1 CB@32_mAd531_2 CB@32_mAd532_1 CB@32_mAd532_2 CB@32_mAd533_1 CB@32_mAd533_2 CB@32_mAd534_1 CB@32_mAd534_2 CB@32_mAd535_1 CB@32_mAd535_2 CB@32_mAd536_1 CB@32_mAd536_2 CB@32_mAd537_1 CB@32_mAd537_2 CB@32_mAd540_1 CB@32_mAd540_2 CB@32_mAd541_1 CB@32_mAd541_2 CB@32_mAd542_1 CB@32_mAd542_2 CB@32_mAd543_1 CB@32_mAd543_2 CB@32_mAd544_1 CB@32_mAd544_2 CB@32_mAd545_1 
+CB@32_mAd545_2 CB@32_mAd546_1 CB@32_mAd546_2 CB@32_mAd547_1 CB@32_mAd547_2 CB@32_mAd550_1 CB@32_mAd550_2 CB@32_mAd551_1 CB@32_mAd551_2 CB@32_mAd552_1 CB@32_mAd552_2 CB@32_mAd553_1 CB@32_mAd553_2 CB@32_mAd554_1 CB@32_mAd554_2 CB@32_mAd555_1 CB@32_mAd555_2 CB@32_mAd556_1 CB@32_mAd556_2 CB@32_mAd557_1 CB@32_mAd557_2 CB@32_mAd560_1 CB@32_mAd560_2 CB@32_mAd561_1 CB@32_mAd561_2 CB@32_mAd562_1 CB@32_mAd562_2 CB@32_mAd563_1 CB@32_mAd563_2 CB@32_mAd564_1 CB@32_mAd564_2 CB@32_mAd565_1 CB@32_mAd565_2 CB@32_mAd566_1 
+CB@32_mAd566_2 CB@32_mAd567_1 CB@32_mAd567_2 CB@32_mAd570_1 CB@32_mAd570_2 CB@32_mAd571_1 CB@32_mAd571_2 CB@32_mAd572_1 CB@32_mAd572_2 CB@32_mAd573_1 CB@32_mAd573_2 CB@32_mAd575_1 CB@32_mAd575_2 CB@32_mAd576_1 CB@32_mAd576_2 CB@32_mAd577_1 CB@32_mAd577_2 CB@32_mAd600_1 CB@32_mAd600_2 CB@32_mAd601_1 CB@32_mAd601_2 CB@32_mAd602_1 CB@32_mAd602_2 CB@32_mAd604_1 CB@32_mAd604_2 CB@32_mAd605_1 CB@32_mAd605_2 CB@32_mAd606_1 CB@32_mAd606_2 CB@32_mAd607_1 CB@32_mAd607_2 CB@32_mAd610_1 CB@32_mAd610_2 CB@32_mAd611_1 
+CB@32_mAd611_2 CB@32_mAd612_1 CB@32_mAd612_2 CB@32_mAd613_1 CB@32_mAd613_2 CB@32_mAd614_1 CB@32_mAd614_2 CB@32_mAd615_1 CB@32_mAd615_2 CB@32_mAd616_1 CB@32_mAd616_2 CB@32_mAd617_1 CB@32_mAd617_2 CB@32_mAd620_1 CB@32_mAd620_2 CB@32_mAd621_1 CB@32_mAd621_2 CB@32_mAd622_1 CB@32_mAd622_2 CB@32_mAd623_1 CB@32_mAd623_2 CB@32_mAd624_1 CB@32_mAd624_2 CB@32_mAd625_1 CB@32_mAd625_2 CB@32_mAd626_1 CB@32_mAd626_2 CB@32_mAd627_1 CB@32_mAd627_2 CB@32_mAd630_1 CB@32_mAd630_2 CB@32_mAd631_1 CB@32_mAd631_2 CB@32_mAd632_1 
+CB@32_mAd632_2 CB@32_mAd633_1 CB@32_mAd633_2 CB@32_mAd634_1 CB@32_mAd634_2 CB@32_mAd635_1 CB@32_mAd635_2 CB@32_mAd636_1 CB@32_mAd636_2 CB@32_mAd637_1 CB@32_mAd637_2 CB@32_mAd640_1 CB@32_mAd640_2 CB@32_mAd641_1 CB@32_mAd641_2 CB@32_mAd642_1 CB@32_mAd642_2 CB@32_mAd643_1 CB@32_mAd643_2 CB@32_mAd644_1 CB@32_mAd644_2 CB@32_mAd645_1 CB@32_mAd645_2 CB@32_mAd646_1 CB@32_mAd646_2 CB@32_mAd647_1 CB@32_mAd647_2 CB@32_mAd650_1 CB@32_mAd650_2 CB@32_mAd651_1 CB@32_mAd651_2 CB@32_mAd652_1 CB@32_mAd652_2 CB@32_mAd653_1 
+CB@32_mAd653_2 CB@32_mAd654_1 CB@32_mAd654_2 CB@32_mAd655_1 CB@32_mAd655_2 CB@32_mAd656_1 CB@32_mAd656_2 CB@32_mAd657_1 CB@32_mAd657_2 CB@32_mAd660_1 CB@32_mAd660_2 CB@32_mAd661_1 CB@32_mAd661_2 CB@32_mAd662_1 CB@32_mAd662_2 CB@32_mAd663_1 CB@32_mAd663_2 CB@32_mAd664_1 CB@32_mAd664_2 CB@32_mAd665_1 CB@32_mAd665_2 CB@32_mAd666_1 CB@32_mAd666_2 CB@32_mAd667_1 CB@32_mAd667_2 CB@32_mAd675_1 CB@32_mAd675_2 CB@32_mAd676_1 CB@32_mAd676_2 CB@32_mAd677_1 CB@32_mAd677_2 CB@32_mAd700_1 CB@32_mAd700_2 CB@32_mAd710_1 
+CB@32_mAd710_2 CB@32_mAd711_1 CB@32_mAd711_2 CB@32_mAd717_1 CB@32_mAd717_2 CB@32_mAd720_1 CB@32_mAd720_2 CB@32_mAd721_1 CB@32_mAd721_2 CB@32_mAd722_1 CB@32_mAd722_2 CB@32_mAd723_1 CB@32_mAd723_2 CB@32_mAd724_1 CB@32_mAd724_2 CB@32_mAd725_1 CB@32_mAd725_2 CB@32_mAd726_1 CB@32_mAd726_2 CB@32_mAd727_1 CB@32_mAd727_2 CB@32_mAd730_1 CB@32_mAd730_2 CB@32_mAd731_1 CB@32_mAd731_2 CB@32_mAd732_1 CB@32_mAd732_2 CB@32_mAd733_1 CB@32_mAd733_2 CB@32_mAd734_1 CB@32_mAd734_2 CB@32_mAd735_1 CB@32_mAd735_2 CB@32_mAd736_1 
+CB@32_mAd736_2 CB@32_mAd737_1 CB@32_mAd737_2 CB@32_mAd740_1 CB@32_mAd740_2 CB@32_mAd741_1 CB@32_mAd741_2 CB@32_mAd742_1 CB@32_mAd742_2 CB@32_mAd743_1 CB@32_mAd743_2 CB@32_mAd744_1 CB@32_mAd744_2 CB@32_mAd745_1 CB@32_mAd745_2 CB@32_mAd746_1 CB@32_mAd746_2 CB@32_mAd747_1 CB@32_mAd747_2 CB@32_mAd750_1 CB@32_mAd750_2 CB@32_mAd751_1 CB@32_mAd751_2 CB@32_mAd752_1 CB@32_mAd752_2 CB@32_mAd753_1 CB@32_mAd753_2 CB@32_mAd754_1 CB@32_mAd754_2 CB@32_mAd755_1 CB@32_mAd755_2 CB@32_mAd756_1 CB@32_mAd756_2 CB@32_mAd757_1 
+CB@32_mAd757_2 CB@32_mAd760_1 CB@32_mAd760_2 CB@32_mAd761_1 CB@32_mAd761_2 CB@32_mAd762_1 CB@32_mAd762_2 CB@32_mAd763_1 CB@32_mAd763_2 CB@32_mAd764_1 CB@32_mAd764_2 CB@32_mAd765_1 CB@32_mAd765_2 CB@32_mAd766_1 CB@32_mAd766_2 CB@32_mAd767_1 CB@32_mAd767_2 CB@32_mAd771_1 CB@32_mAd771_2 CB@32_mAd772_1 CB@32_mAd772_2 CB@32_mAd773_1 CB@32_mAd773_2 CB@32_mAd774_1 CB@32_mAd774_2 CB@32_mAd775_1 CB@32_mAd775_2 CB@32_mAd776_1 CB@32_mAd776_2 CB@32_mAd777_1 CB@32_mAd777_2 CB@32_X0 CB@32_X1 CB@32_X10 CB@32_X11 
+CB@32_X12 CB@32_X13 CB@32_X2 CB@32_X3 CB@32_X4 CB@32_X5 CB@32_X6 CB@32_X7 CB@32_X8 CB@32_X9 CB@32_Y1 CB@32_Y10 CB@32_Y11 CB@32_Y12 CB@32_Y2 CB@32_Y3 CB@32_Y4 CB@32_Y5 CB@32_Y6 CB@32_Y7 CB@32_Y8 CB@32_Y9 CB@32_Z1 CB@32_Z10 CB@32_Z11 CB@32_Z12 CB@32_Z2 CB@32_Z3 CB@32_Z4 CB@32_Z5 CB@32_Z6 CB@32_Z7 CB@32_Z8 CB@32_Z9 _5400TP094__CB
XCB@33 CB@33_K0 CB@33_K1 CB@33_K10 CB@33_K11 CB@33_K12 CB@33_K13 CB@33_K2 CB@33_K3 CB@33_K4 CB@33_K5 CB@33_K6 CB@33_K7 CB@33_K8 CB@33_K9 CB@33_mAd000_1 CB@33_mAd000_2 CB@33_mAd001_1 CB@33_mAd001_2 CB@33_mAd002_1 CB@33_mAd002_2 CB@33_mAd003_1 CB@33_mAd003_2 CB@33_mAd004_1 CB@33_mAd004_2 CB@33_mAd005_1 CB@33_mAd005_2 CB@33_mAd006_1 CB@33_mAd006_2 CB@33_mAd007_1 CB@33_mAd007_2 CB@33_mAd010_1 CB@33_mAd010_2 CB@33_mAd011_1 CB@33_mAd011_2 CB@33_mAd012_1 CB@33_mAd012_2 CB@33_mAd013_1 CB@33_mAd013_2 CB@33_mAd014_1 
+CB@33_mAd014_2 CB@33_mAd015_1 CB@33_mAd015_2 CB@33_mAd016_1 CB@33_mAd016_2 CB@33_mAd017_1 CB@33_mAd017_2 CB@33_mAd020_1 CB@33_mAd020_2 CB@33_mAd021_1 CB@33_mAd021_2 CB@33_mAd022_1 CB@33_mAd022_2 CB@33_mAd023_1 CB@33_mAd023_2 CB@33_mAd024_1 CB@33_mAd024_2 CB@33_mAd025_1 CB@33_mAd025_2 CB@33_mAd026_1 CB@33_mAd026_2 CB@33_mAd027_1 CB@33_mAd027_2 CB@33_mAd030_1 CB@33_mAd030_2 CB@33_mAd031_1 CB@33_mAd031_2 CB@33_mAd032_1 CB@33_mAd032_2 CB@33_mAd033_1 CB@33_mAd033_2 CB@33_mAd034_1 CB@33_mAd034_2 CB@33_mAd035_1 
+CB@33_mAd035_2 CB@33_mAd036_1 CB@33_mAd036_2 CB@33_mAd037_1 CB@33_mAd037_2 CB@33_mAd040_1 CB@33_mAd040_2 CB@33_mAd041_1 CB@33_mAd041_2 CB@33_mAd042_1 CB@33_mAd042_2 CB@33_mAd043_1 CB@33_mAd043_2 CB@33_mAd044_1 CB@33_mAd044_2 CB@33_mAd045_1 CB@33_mAd045_2 CB@33_mAd046_1 CB@33_mAd046_2 CB@33_mAd047_1 CB@33_mAd047_2 CB@33_mAd050_1 CB@33_mAd050_2 CB@33_mAd051_1 CB@33_mAd051_2 CB@33_mAd052_1 CB@33_mAd052_2 CB@33_mAd053_1 CB@33_mAd053_2 CB@33_mAd054_1 CB@33_mAd054_2 CB@33_mAd055_1 CB@33_mAd055_2 CB@33_mAd056_1 
+CB@33_mAd056_2 CB@33_mAd057_1 CB@33_mAd057_2 CB@33_mAd060_1 CB@33_mAd060_2 CB@33_mAd066_1 CB@33_mAd066_2 CB@33_mAd067_1 CB@33_mAd067_2 CB@33_mAd100_1 CB@33_mAd100_2 CB@33_mAd101_1 CB@33_mAd101_2 CB@33_mAd102_1 CB@33_mAd102_2 CB@33_mAd110_1 CB@33_mAd110_2 CB@33_mAd111_1 CB@33_mAd111_2 CB@33_mAd112_1 CB@33_mAd112_2 CB@33_mAd113_1 CB@33_mAd113_2 CB@33_mAd114_1 CB@33_mAd114_2 CB@33_mAd115_1 CB@33_mAd115_2 CB@33_mAd116_1 CB@33_mAd116_2 CB@33_mAd117_1 CB@33_mAd117_2 CB@33_mAd120_1 CB@33_mAd120_2 CB@33_mAd121_1 
+CB@33_mAd121_2 CB@33_mAd122_1 CB@33_mAd122_2 CB@33_mAd123_1 CB@33_mAd123_2 CB@33_mAd124_1 CB@33_mAd124_2 CB@33_mAd125_1 CB@33_mAd125_2 CB@33_mAd126_1 CB@33_mAd126_2 CB@33_mAd127_1 CB@33_mAd127_2 CB@33_mAd130_1 CB@33_mAd130_2 CB@33_mAd131_1 CB@33_mAd131_2 CB@33_mAd132_1 CB@33_mAd132_2 CB@33_mAd133_1 CB@33_mAd133_2 CB@33_mAd134_1 CB@33_mAd134_2 CB@33_mAd135_1 CB@33_mAd135_2 CB@33_mAd136_1 CB@33_mAd136_2 CB@33_mAd137_1 CB@33_mAd137_2 CB@33_mAd140_1 CB@33_mAd140_2 CB@33_mAd141_1 CB@33_mAd141_2 CB@33_mAd142_1 
+CB@33_mAd142_2 CB@33_mAd143_1 CB@33_mAd143_2 CB@33_mAd144_1 CB@33_mAd144_2 CB@33_mAd145_1 CB@33_mAd145_2 CB@33_mAd146_1 CB@33_mAd146_2 CB@33_mAd147_1 CB@33_mAd147_2 CB@33_mAd150_1 CB@33_mAd150_2 CB@33_mAd151_1 CB@33_mAd151_2 CB@33_mAd152_1 CB@33_mAd152_2 CB@33_mAd153_1 CB@33_mAd153_2 CB@33_mAd154_1 CB@33_mAd154_2 CB@33_mAd155_1 CB@33_mAd155_2 CB@33_mAd156_1 CB@33_mAd156_2 CB@33_mAd157_1 CB@33_mAd157_2 CB@33_mAd160_1 CB@33_mAd160_2 CB@33_mAd161_1 CB@33_mAd161_2 CB@33_mAd162_1 CB@33_mAd162_2 CB@33_mAd163_1 
+CB@33_mAd163_2 CB@33_mAd164_1 CB@33_mAd164_2 CB@33_mAd165_1 CB@33_mAd165_2 CB@33_mAd166_1 CB@33_mAd166_2 CB@33_mAd167_1 CB@33_mAd167_2 CB@33_mAd170_1 CB@33_mAd170_2 CB@33_mAd171_1 CB@33_mAd171_2 CB@33_mAd172_1 CB@33_mAd172_2 CB@33_mAd173_1 CB@33_mAd173_2 CB@33_mAd175_1 CB@33_mAd175_2 CB@33_mAd176_1 CB@33_mAd176_2 CB@33_mAd177_1 CB@33_mAd177_2 CB@33_mAd200_1 CB@33_mAd200_2 CB@33_mAd201_1 CB@33_mAd201_2 CB@33_mAd202_1 CB@33_mAd202_2 CB@33_mAd204_1 CB@33_mAd204_2 CB@33_mAd205_1 CB@33_mAd205_2 CB@33_mAd206_1 
+CB@33_mAd206_2 CB@33_mAd207_1 CB@33_mAd207_2 CB@33_mAd210_1 CB@33_mAd210_2 CB@33_mAd211_1 CB@33_mAd211_2 CB@33_mAd212_1 CB@33_mAd212_2 CB@33_mAd213_1 CB@33_mAd213_2 CB@33_mAd214_1 CB@33_mAd214_2 CB@33_mAd215_1 CB@33_mAd215_2 CB@33_mAd216_1 CB@33_mAd216_2 CB@33_mAd217_1 CB@33_mAd217_2 CB@33_mAd220_1 CB@33_mAd220_2 CB@33_mAd221_1 CB@33_mAd221_2 CB@33_mAd222_1 CB@33_mAd222_2 CB@33_mAd223_1 CB@33_mAd223_2 CB@33_mAd224_1 CB@33_mAd224_2 CB@33_mAd225_1 CB@33_mAd225_2 CB@33_mAd226_1 CB@33_mAd226_2 CB@33_mAd227_1 
+CB@33_mAd227_2 CB@33_mAd230_1 CB@33_mAd230_2 CB@33_mAd231_1 CB@33_mAd231_2 CB@33_mAd232_1 CB@33_mAd232_2 CB@33_mAd233_1 CB@33_mAd233_2 CB@33_mAd234_1 CB@33_mAd234_2 CB@33_mAd235_1 CB@33_mAd235_2 CB@33_mAd236_1 CB@33_mAd236_2 CB@33_mAd237_1 CB@33_mAd237_2 CB@33_mAd240_1 CB@33_mAd240_2 CB@33_mAd241_1 CB@33_mAd241_2 CB@33_mAd242_1 CB@33_mAd242_2 CB@33_mAd243_1 CB@33_mAd243_2 CB@33_mAd244_1 CB@33_mAd244_2 CB@33_mAd245_1 CB@33_mAd245_2 CB@33_mAd246_1 CB@33_mAd246_2 CB@33_mAd247_1 CB@33_mAd247_2 CB@33_mAd250_1 
+CB@33_mAd250_2 CB@33_mAd251_1 CB@33_mAd251_2 CB@33_mAd252_1 CB@33_mAd252_2 CB@33_mAd253_1 CB@33_mAd253_2 CB@33_mAd254_1 CB@33_mAd254_2 CB@33_mAd255_1 CB@33_mAd255_2 CB@33_mAd256_1 CB@33_mAd256_2 CB@33_mAd257_1 CB@33_mAd257_2 CB@33_mAd260_1 CB@33_mAd260_2 CB@33_mAd261_1 CB@33_mAd261_2 CB@33_mAd262_1 CB@33_mAd262_2 CB@33_mAd263_1 CB@33_mAd263_2 CB@33_mAd264_1 CB@33_mAd264_2 CB@33_mAd265_1 CB@33_mAd265_2 CB@33_mAd266_1 CB@33_mAd266_2 CB@33_mAd267_1 CB@33_mAd267_2 CB@33_mAd275_1 CB@33_mAd275_2 CB@33_mAd276_1 
+CB@33_mAd276_2 CB@33_mAd277_1 CB@33_mAd277_2 CB@33_mAd300_1 CB@33_mAd300_2 CB@33_mAd310_1 CB@33_mAd310_2 CB@33_mAd311_1 CB@33_mAd311_2 CB@33_mAd317_1 CB@33_mAd317_2 CB@33_mAd320_1 CB@33_mAd320_2 CB@33_mAd321_1 CB@33_mAd321_2 CB@33_mAd322_1 CB@33_mAd322_2 CB@33_mAd323_1 CB@33_mAd323_2 CB@33_mAd324_1 CB@33_mAd324_2 CB@33_mAd325_1 CB@33_mAd325_2 CB@33_mAd326_1 CB@33_mAd326_2 CB@33_mAd327_1 CB@33_mAd327_2 CB@33_mAd330_1 CB@33_mAd330_2 CB@33_mAd331_1 CB@33_mAd331_2 CB@33_mAd332_1 CB@33_mAd332_2 CB@33_mAd333_1 
+CB@33_mAd333_2 CB@33_mAd334_1 CB@33_mAd334_2 CB@33_mAd335_1 CB@33_mAd335_2 CB@33_mAd336_1 CB@33_mAd336_2 CB@33_mAd337_1 CB@33_mAd337_2 CB@33_mAd340_1 CB@33_mAd340_2 CB@33_mAd341_1 CB@33_mAd341_2 CB@33_mAd342_1 CB@33_mAd342_2 CB@33_mAd343_1 CB@33_mAd343_2 CB@33_mAd344_1 CB@33_mAd344_2 CB@33_mAd345_1 CB@33_mAd345_2 CB@33_mAd346_1 CB@33_mAd346_2 CB@33_mAd347_1 CB@33_mAd347_2 CB@33_mAd350_1 CB@33_mAd350_2 CB@33_mAd351_1 CB@33_mAd351_2 CB@33_mAd352_1 CB@33_mAd352_2 CB@33_mAd353_1 CB@33_mAd353_2 CB@33_mAd354_1 
+CB@33_mAd354_2 CB@33_mAd355_1 CB@33_mAd355_2 CB@33_mAd356_1 CB@33_mAd356_2 CB@33_mAd357_1 CB@33_mAd357_2 CB@33_mAd360_1 CB@33_mAd360_2 CB@33_mAd361_1 CB@33_mAd361_2 CB@33_mAd362_1 CB@33_mAd362_2 CB@33_mAd363_1 CB@33_mAd363_2 CB@33_mAd364_1 CB@33_mAd364_2 CB@33_mAd365_1 CB@33_mAd365_2 CB@33_mAd366_1 CB@33_mAd366_2 CB@33_mAd367_1 CB@33_mAd367_2 CB@33_mAd371_1 CB@33_mAd371_2 CB@33_mAd372_1 CB@33_mAd372_2 CB@33_mAd373_1 CB@33_mAd373_2 CB@33_mAd374_1 CB@33_mAd374_2 CB@33_mAd375_1 CB@33_mAd375_2 CB@33_mAd376_1 
+CB@33_mAd376_2 CB@33_mAd377_1 CB@33_mAd377_2 CB@33_mAd400_1 CB@33_mAd400_2 CB@33_mAd401_1 CB@33_mAd401_2 CB@33_mAd402_1 CB@33_mAd402_2 CB@33_mAd403_1 CB@33_mAd403_2 CB@33_mAd404_1 CB@33_mAd404_2 CB@33_mAd405_1 CB@33_mAd405_2 CB@33_mAd406_1 CB@33_mAd406_2 CB@33_mAd407_1 CB@33_mAd407_2 CB@33_mAd410_1 CB@33_mAd410_2 CB@33_mAd411_1 CB@33_mAd411_2 CB@33_mAd412_1 CB@33_mAd412_2 CB@33_mAd413_1 CB@33_mAd413_2 CB@33_mAd414_1 CB@33_mAd414_2 CB@33_mAd415_1 CB@33_mAd415_2 CB@33_mAd416_1 CB@33_mAd416_2 CB@33_mAd417_1 
+CB@33_mAd417_2 CB@33_mAd420_1 CB@33_mAd420_2 CB@33_mAd421_1 CB@33_mAd421_2 CB@33_mAd422_1 CB@33_mAd422_2 CB@33_mAd423_1 CB@33_mAd423_2 CB@33_mAd424_1 CB@33_mAd424_2 CB@33_mAd425_1 CB@33_mAd425_2 CB@33_mAd426_1 CB@33_mAd426_2 CB@33_mAd427_1 CB@33_mAd427_2 CB@33_mAd430_1 CB@33_mAd430_2 CB@33_mAd431_1 CB@33_mAd431_2 CB@33_mAd432_1 CB@33_mAd432_2 CB@33_mAd433_1 CB@33_mAd433_2 CB@33_mAd434_1 CB@33_mAd434_2 CB@33_mAd435_1 CB@33_mAd435_2 CB@33_mAd436_1 CB@33_mAd436_2 CB@33_mAd437_1 CB@33_mAd437_2 CB@33_mAd440_1 
+CB@33_mAd440_2 CB@33_mAd441_1 CB@33_mAd441_2 CB@33_mAd442_1 CB@33_mAd442_2 CB@33_mAd443_1 CB@33_mAd443_2 CB@33_mAd444_1 CB@33_mAd444_2 CB@33_mAd445_1 CB@33_mAd445_2 CB@33_mAd446_1 CB@33_mAd446_2 CB@33_mAd447_1 CB@33_mAd447_2 CB@33_mAd450_1 CB@33_mAd450_2 CB@33_mAd451_1 CB@33_mAd451_2 CB@33_mAd452_1 CB@33_mAd452_2 CB@33_mAd453_1 CB@33_mAd453_2 CB@33_mAd454_1 CB@33_mAd454_2 CB@33_mAd455_1 CB@33_mAd455_2 CB@33_mAd456_1 CB@33_mAd456_2 CB@33_mAd457_1 CB@33_mAd457_2 CB@33_mAd460_1 CB@33_mAd460_2 CB@33_mAd466_1 
+CB@33_mAd466_2 CB@33_mAd467_1 CB@33_mAd467_2 CB@33_mAd500_1 CB@33_mAd500_2 CB@33_mAd501_1 CB@33_mAd501_2 CB@33_mAd502_1 CB@33_mAd502_2 CB@33_mAd508_1 CB@33_mAd508_2 CB@33_mAd509_1 CB@33_mAd509_2 CB@33_mAd512_1 CB@33_mAd512_2 CB@33_mAd513_1 CB@33_mAd513_2 CB@33_mAd514_1 CB@33_mAd514_2 CB@33_mAd515_1 CB@33_mAd515_2 CB@33_mAd516_1 CB@33_mAd516_2 CB@33_mAd517_1 CB@33_mAd517_2 CB@33_mAd520_1 CB@33_mAd520_2 CB@33_mAd521_1 CB@33_mAd521_2 CB@33_mAd522_1 CB@33_mAd522_2 CB@33_mAd523_1 CB@33_mAd523_2 CB@33_mAd524_1 
+CB@33_mAd524_2 CB@33_mAd525_1 CB@33_mAd525_2 CB@33_mAd526_1 CB@33_mAd526_2 CB@33_mAd527_1 CB@33_mAd527_2 CB@33_mAd530_1 CB@33_mAd530_2 CB@33_mAd531_1 CB@33_mAd531_2 CB@33_mAd532_1 CB@33_mAd532_2 CB@33_mAd533_1 CB@33_mAd533_2 CB@33_mAd534_1 CB@33_mAd534_2 CB@33_mAd535_1 CB@33_mAd535_2 CB@33_mAd536_1 CB@33_mAd536_2 CB@33_mAd537_1 CB@33_mAd537_2 CB@33_mAd540_1 CB@33_mAd540_2 CB@33_mAd541_1 CB@33_mAd541_2 CB@33_mAd542_1 CB@33_mAd542_2 CB@33_mAd543_1 CB@33_mAd543_2 CB@33_mAd544_1 CB@33_mAd544_2 CB@33_mAd545_1 
+CB@33_mAd545_2 CB@33_mAd546_1 CB@33_mAd546_2 CB@33_mAd547_1 CB@33_mAd547_2 CB@33_mAd550_1 CB@33_mAd550_2 CB@33_mAd551_1 CB@33_mAd551_2 CB@33_mAd552_1 CB@33_mAd552_2 CB@33_mAd553_1 CB@33_mAd553_2 CB@33_mAd554_1 CB@33_mAd554_2 CB@33_mAd555_1 CB@33_mAd555_2 CB@33_mAd556_1 CB@33_mAd556_2 CB@33_mAd557_1 CB@33_mAd557_2 CB@33_mAd560_1 CB@33_mAd560_2 CB@33_mAd561_1 CB@33_mAd561_2 CB@33_mAd562_1 CB@33_mAd562_2 CB@33_mAd563_1 CB@33_mAd563_2 CB@33_mAd564_1 CB@33_mAd564_2 CB@33_mAd565_1 CB@33_mAd565_2 CB@33_mAd566_1 
+CB@33_mAd566_2 CB@33_mAd567_1 CB@33_mAd567_2 CB@33_mAd570_1 CB@33_mAd570_2 CB@33_mAd571_1 CB@33_mAd571_2 CB@33_mAd572_1 CB@33_mAd572_2 CB@33_mAd573_1 CB@33_mAd573_2 CB@33_mAd575_1 CB@33_mAd575_2 CB@33_mAd576_1 CB@33_mAd576_2 CB@33_mAd577_1 CB@33_mAd577_2 CB@33_mAd600_1 CB@33_mAd600_2 CB@33_mAd601_1 CB@33_mAd601_2 CB@33_mAd602_1 CB@33_mAd602_2 CB@33_mAd604_1 CB@33_mAd604_2 CB@33_mAd605_1 CB@33_mAd605_2 CB@33_mAd606_1 CB@33_mAd606_2 CB@33_mAd607_1 CB@33_mAd607_2 CB@33_mAd610_1 CB@33_mAd610_2 CB@33_mAd611_1 
+CB@33_mAd611_2 CB@33_mAd612_1 CB@33_mAd612_2 CB@33_mAd613_1 CB@33_mAd613_2 CB@33_mAd614_1 CB@33_mAd614_2 CB@33_mAd615_1 CB@33_mAd615_2 CB@33_mAd616_1 CB@33_mAd616_2 CB@33_mAd617_1 CB@33_mAd617_2 CB@33_mAd620_1 CB@33_mAd620_2 CB@33_mAd621_1 CB@33_mAd621_2 CB@33_mAd622_1 CB@33_mAd622_2 CB@33_mAd623_1 CB@33_mAd623_2 CB@33_mAd624_1 CB@33_mAd624_2 CB@33_mAd625_1 CB@33_mAd625_2 CB@33_mAd626_1 CB@33_mAd626_2 CB@33_mAd627_1 CB@33_mAd627_2 CB@33_mAd630_1 CB@33_mAd630_2 CB@33_mAd631_1 CB@33_mAd631_2 CB@33_mAd632_1 
+CB@33_mAd632_2 CB@33_mAd633_1 CB@33_mAd633_2 CB@33_mAd634_1 CB@33_mAd634_2 CB@33_mAd635_1 CB@33_mAd635_2 CB@33_mAd636_1 CB@33_mAd636_2 CB@33_mAd637_1 CB@33_mAd637_2 CB@33_mAd640_1 CB@33_mAd640_2 CB@33_mAd641_1 CB@33_mAd641_2 CB@33_mAd642_1 CB@33_mAd642_2 CB@33_mAd643_1 CB@33_mAd643_2 CB@33_mAd644_1 CB@33_mAd644_2 CB@33_mAd645_1 CB@33_mAd645_2 CB@33_mAd646_1 CB@33_mAd646_2 CB@33_mAd647_1 CB@33_mAd647_2 CB@33_mAd650_1 CB@33_mAd650_2 CB@33_mAd651_1 CB@33_mAd651_2 CB@33_mAd652_1 CB@33_mAd652_2 CB@33_mAd653_1 
+CB@33_mAd653_2 CB@33_mAd654_1 CB@33_mAd654_2 CB@33_mAd655_1 CB@33_mAd655_2 CB@33_mAd656_1 CB@33_mAd656_2 CB@33_mAd657_1 CB@33_mAd657_2 CB@33_mAd660_1 CB@33_mAd660_2 CB@33_mAd661_1 CB@33_mAd661_2 CB@33_mAd662_1 CB@33_mAd662_2 CB@33_mAd663_1 CB@33_mAd663_2 CB@33_mAd664_1 CB@33_mAd664_2 CB@33_mAd665_1 CB@33_mAd665_2 CB@33_mAd666_1 CB@33_mAd666_2 CB@33_mAd667_1 CB@33_mAd667_2 CB@33_mAd675_1 CB@33_mAd675_2 CB@33_mAd676_1 CB@33_mAd676_2 CB@33_mAd677_1 CB@33_mAd677_2 CB@33_mAd700_1 CB@33_mAd700_2 CB@33_mAd710_1 
+CB@33_mAd710_2 CB@33_mAd711_1 CB@33_mAd711_2 CB@33_mAd717_1 CB@33_mAd717_2 CB@33_mAd720_1 CB@33_mAd720_2 CB@33_mAd721_1 CB@33_mAd721_2 CB@33_mAd722_1 CB@33_mAd722_2 CB@33_mAd723_1 CB@33_mAd723_2 CB@33_mAd724_1 CB@33_mAd724_2 CB@33_mAd725_1 CB@33_mAd725_2 CB@33_mAd726_1 CB@33_mAd726_2 CB@33_mAd727_1 CB@33_mAd727_2 CB@33_mAd730_1 CB@33_mAd730_2 CB@33_mAd731_1 CB@33_mAd731_2 CB@33_mAd732_1 CB@33_mAd732_2 CB@33_mAd733_1 CB@33_mAd733_2 CB@33_mAd734_1 CB@33_mAd734_2 CB@33_mAd735_1 CB@33_mAd735_2 CB@33_mAd736_1 
+CB@33_mAd736_2 CB@33_mAd737_1 CB@33_mAd737_2 CB@33_mAd740_1 CB@33_mAd740_2 CB@33_mAd741_1 CB@33_mAd741_2 CB@33_mAd742_1 CB@33_mAd742_2 CB@33_mAd743_1 CB@33_mAd743_2 CB@33_mAd744_1 CB@33_mAd744_2 CB@33_mAd745_1 CB@33_mAd745_2 CB@33_mAd746_1 CB@33_mAd746_2 CB@33_mAd747_1 CB@33_mAd747_2 CB@33_mAd750_1 CB@33_mAd750_2 CB@33_mAd751_1 CB@33_mAd751_2 CB@33_mAd752_1 CB@33_mAd752_2 CB@33_mAd753_1 CB@33_mAd753_2 CB@33_mAd754_1 CB@33_mAd754_2 CB@33_mAd755_1 CB@33_mAd755_2 CB@33_mAd756_1 CB@33_mAd756_2 CB@33_mAd757_1 
+CB@33_mAd757_2 CB@33_mAd760_1 CB@33_mAd760_2 CB@33_mAd761_1 CB@33_mAd761_2 CB@33_mAd762_1 CB@33_mAd762_2 CB@33_mAd763_1 CB@33_mAd763_2 CB@33_mAd764_1 CB@33_mAd764_2 CB@33_mAd765_1 CB@33_mAd765_2 CB@33_mAd766_1 CB@33_mAd766_2 CB@33_mAd767_1 CB@33_mAd767_2 CB@33_mAd771_1 CB@33_mAd771_2 CB@33_mAd772_1 CB@33_mAd772_2 CB@33_mAd773_1 CB@33_mAd773_2 CB@33_mAd774_1 CB@33_mAd774_2 CB@33_mAd775_1 CB@33_mAd775_2 CB@33_mAd776_1 CB@33_mAd776_2 CB@33_mAd777_1 CB@33_mAd777_2 CB@33_X0 CB@33_X1 CB@33_X10 CB@33_X11 
+CB@33_X12 CB@33_X13 CB@33_X2 CB@33_X3 CB@33_X4 CB@33_X5 CB@33_X6 CB@33_X7 CB@33_X8 CB@33_X9 CB@33_Y1 CB@33_Y10 CB@33_Y11 CB@33_Y12 CB@33_Y2 CB@33_Y3 CB@33_Y4 CB@33_Y5 CB@33_Y6 CB@33_Y7 CB@33_Y8 CB@33_Y9 CB@33_Z1 CB@33_Z10 CB@33_Z11 CB@33_Z12 CB@33_Z2 CB@33_Z3 CB@33_Z4 CB@33_Z5 CB@33_Z6 CB@33_Z7 CB@33_Z8 CB@33_Z9 _5400TP094__CB
XCB@34 CB@34_K0 CB@34_K1 CB@34_K10 CB@34_K11 CB@34_K12 CB@34_K13 CB@34_K2 CB@34_K3 CB@34_K4 CB@34_K5 CB@34_K6 CB@34_K7 CB@34_K8 CB@34_K9 CB@34_mAd000_1 CB@34_mAd000_2 CB@34_mAd001_1 CB@34_mAd001_2 CB@34_mAd002_1 CB@34_mAd002_2 CB@34_mAd003_1 CB@34_mAd003_2 CB@34_mAd004_1 CB@34_mAd004_2 CB@34_mAd005_1 CB@34_mAd005_2 CB@34_mAd006_1 CB@34_mAd006_2 CB@34_mAd007_1 CB@34_mAd007_2 CB@34_mAd010_1 CB@34_mAd010_2 CB@34_mAd011_1 CB@34_mAd011_2 CB@34_mAd012_1 CB@34_mAd012_2 CB@34_mAd013_1 CB@34_mAd013_2 CB@34_mAd014_1 
+CB@34_mAd014_2 CB@34_mAd015_1 CB@34_mAd015_2 CB@34_mAd016_1 CB@34_mAd016_2 CB@34_mAd017_1 CB@34_mAd017_2 CB@34_mAd020_1 CB@34_mAd020_2 CB@34_mAd021_1 CB@34_mAd021_2 CB@34_mAd022_1 CB@34_mAd022_2 CB@34_mAd023_1 CB@34_mAd023_2 CB@34_mAd024_1 CB@34_mAd024_2 CB@34_mAd025_1 CB@34_mAd025_2 CB@34_mAd026_1 CB@34_mAd026_2 CB@34_mAd027_1 CB@34_mAd027_2 CB@34_mAd030_1 CB@34_mAd030_2 CB@34_mAd031_1 CB@34_mAd031_2 CB@34_mAd032_1 CB@34_mAd032_2 CB@34_mAd033_1 CB@34_mAd033_2 CB@34_mAd034_1 CB@34_mAd034_2 CB@34_mAd035_1 
+CB@34_mAd035_2 CB@34_mAd036_1 CB@34_mAd036_2 CB@34_mAd037_1 CB@34_mAd037_2 CB@34_mAd040_1 CB@34_mAd040_2 CB@34_mAd041_1 CB@34_mAd041_2 CB@34_mAd042_1 CB@34_mAd042_2 CB@34_mAd043_1 CB@34_mAd043_2 CB@34_mAd044_1 CB@34_mAd044_2 CB@34_mAd045_1 CB@34_mAd045_2 CB@34_mAd046_1 CB@34_mAd046_2 CB@34_mAd047_1 CB@34_mAd047_2 CB@34_mAd050_1 CB@34_mAd050_2 CB@34_mAd051_1 CB@34_mAd051_2 CB@34_mAd052_1 CB@34_mAd052_2 CB@34_mAd053_1 CB@34_mAd053_2 CB@34_mAd054_1 CB@34_mAd054_2 CB@34_mAd055_1 CB@34_mAd055_2 CB@34_mAd056_1 
+CB@34_mAd056_2 CB@34_mAd057_1 CB@34_mAd057_2 CB@34_mAd060_1 CB@34_mAd060_2 CB@34_mAd066_1 CB@34_mAd066_2 CB@34_mAd067_1 CB@34_mAd067_2 CB@34_mAd100_1 CB@34_mAd100_2 CB@34_mAd101_1 CB@34_mAd101_2 CB@34_mAd102_1 CB@34_mAd102_2 CB@34_mAd110_1 CB@34_mAd110_2 CB@34_mAd111_1 CB@34_mAd111_2 CB@34_mAd112_1 CB@34_mAd112_2 CB@34_mAd113_1 CB@34_mAd113_2 CB@34_mAd114_1 CB@34_mAd114_2 CB@34_mAd115_1 CB@34_mAd115_2 CB@34_mAd116_1 CB@34_mAd116_2 CB@34_mAd117_1 CB@34_mAd117_2 CB@34_mAd120_1 CB@34_mAd120_2 CB@34_mAd121_1 
+CB@34_mAd121_2 CB@34_mAd122_1 CB@34_mAd122_2 CB@34_mAd123_1 CB@34_mAd123_2 CB@34_mAd124_1 CB@34_mAd124_2 CB@34_mAd125_1 CB@34_mAd125_2 CB@34_mAd126_1 CB@34_mAd126_2 CB@34_mAd127_1 CB@34_mAd127_2 CB@34_mAd130_1 CB@34_mAd130_2 CB@34_mAd131_1 CB@34_mAd131_2 CB@34_mAd132_1 CB@34_mAd132_2 CB@34_mAd133_1 CB@34_mAd133_2 CB@34_mAd134_1 CB@34_mAd134_2 CB@34_mAd135_1 CB@34_mAd135_2 CB@34_mAd136_1 CB@34_mAd136_2 CB@34_mAd137_1 CB@34_mAd137_2 CB@34_mAd140_1 CB@34_mAd140_2 CB@34_mAd141_1 CB@34_mAd141_2 CB@34_mAd142_1 
+CB@34_mAd142_2 CB@34_mAd143_1 CB@34_mAd143_2 CB@34_mAd144_1 CB@34_mAd144_2 CB@34_mAd145_1 CB@34_mAd145_2 CB@34_mAd146_1 CB@34_mAd146_2 CB@34_mAd147_1 CB@34_mAd147_2 CB@34_mAd150_1 CB@34_mAd150_2 CB@34_mAd151_1 CB@34_mAd151_2 CB@34_mAd152_1 CB@34_mAd152_2 CB@34_mAd153_1 CB@34_mAd153_2 CB@34_mAd154_1 CB@34_mAd154_2 CB@34_mAd155_1 CB@34_mAd155_2 CB@34_mAd156_1 CB@34_mAd156_2 CB@34_mAd157_1 CB@34_mAd157_2 CB@34_mAd160_1 CB@34_mAd160_2 CB@34_mAd161_1 CB@34_mAd161_2 CB@34_mAd162_1 CB@34_mAd162_2 CB@34_mAd163_1 
+CB@34_mAd163_2 CB@34_mAd164_1 CB@34_mAd164_2 CB@34_mAd165_1 CB@34_mAd165_2 CB@34_mAd166_1 CB@34_mAd166_2 CB@34_mAd167_1 CB@34_mAd167_2 CB@34_mAd170_1 CB@34_mAd170_2 CB@34_mAd171_1 CB@34_mAd171_2 CB@34_mAd172_1 CB@34_mAd172_2 CB@34_mAd173_1 CB@34_mAd173_2 CB@34_mAd175_1 CB@34_mAd175_2 CB@34_mAd176_1 CB@34_mAd176_2 CB@34_mAd177_1 CB@34_mAd177_2 CB@34_mAd200_1 CB@34_mAd200_2 CB@34_mAd201_1 CB@34_mAd201_2 CB@34_mAd202_1 CB@34_mAd202_2 CB@34_mAd204_1 CB@34_mAd204_2 CB@34_mAd205_1 CB@34_mAd205_2 CB@34_mAd206_1 
+CB@34_mAd206_2 CB@34_mAd207_1 CB@34_mAd207_2 CB@34_mAd210_1 CB@34_mAd210_2 CB@34_mAd211_1 CB@34_mAd211_2 CB@34_mAd212_1 CB@34_mAd212_2 CB@34_mAd213_1 CB@34_mAd213_2 CB@34_mAd214_1 CB@34_mAd214_2 CB@34_mAd215_1 CB@34_mAd215_2 CB@34_mAd216_1 CB@34_mAd216_2 CB@34_mAd217_1 CB@34_mAd217_2 CB@34_mAd220_1 CB@34_mAd220_2 CB@34_mAd221_1 CB@34_mAd221_2 CB@34_mAd222_1 CB@34_mAd222_2 CB@34_mAd223_1 CB@34_mAd223_2 CB@34_mAd224_1 CB@34_mAd224_2 CB@34_mAd225_1 CB@34_mAd225_2 CB@34_mAd226_1 CB@34_mAd226_2 CB@34_mAd227_1 
+CB@34_mAd227_2 CB@34_mAd230_1 CB@34_mAd230_2 CB@34_mAd231_1 CB@34_mAd231_2 CB@34_mAd232_1 CB@34_mAd232_2 CB@34_mAd233_1 CB@34_mAd233_2 CB@34_mAd234_1 CB@34_mAd234_2 CB@34_mAd235_1 CB@34_mAd235_2 CB@34_mAd236_1 CB@34_mAd236_2 CB@34_mAd237_1 CB@34_mAd237_2 CB@34_mAd240_1 CB@34_mAd240_2 CB@34_mAd241_1 CB@34_mAd241_2 CB@34_mAd242_1 CB@34_mAd242_2 CB@34_mAd243_1 CB@34_mAd243_2 CB@34_mAd244_1 CB@34_mAd244_2 CB@34_mAd245_1 CB@34_mAd245_2 CB@34_mAd246_1 CB@34_mAd246_2 CB@34_mAd247_1 CB@34_mAd247_2 CB@34_mAd250_1 
+CB@34_mAd250_2 CB@34_mAd251_1 CB@34_mAd251_2 CB@34_mAd252_1 CB@34_mAd252_2 CB@34_mAd253_1 CB@34_mAd253_2 CB@34_mAd254_1 CB@34_mAd254_2 CB@34_mAd255_1 CB@34_mAd255_2 CB@34_mAd256_1 CB@34_mAd256_2 CB@34_mAd257_1 CB@34_mAd257_2 CB@34_mAd260_1 CB@34_mAd260_2 CB@34_mAd261_1 CB@34_mAd261_2 CB@34_mAd262_1 CB@34_mAd262_2 CB@34_mAd263_1 CB@34_mAd263_2 CB@34_mAd264_1 CB@34_mAd264_2 CB@34_mAd265_1 CB@34_mAd265_2 CB@34_mAd266_1 CB@34_mAd266_2 CB@34_mAd267_1 CB@34_mAd267_2 CB@34_mAd275_1 CB@34_mAd275_2 CB@34_mAd276_1 
+CB@34_mAd276_2 CB@34_mAd277_1 CB@34_mAd277_2 CB@34_mAd300_1 CB@34_mAd300_2 CB@34_mAd310_1 CB@34_mAd310_2 CB@34_mAd311_1 CB@34_mAd311_2 CB@34_mAd317_1 CB@34_mAd317_2 CB@34_mAd320_1 CB@34_mAd320_2 CB@34_mAd321_1 CB@34_mAd321_2 CB@34_mAd322_1 CB@34_mAd322_2 CB@34_mAd323_1 CB@34_mAd323_2 CB@34_mAd324_1 CB@34_mAd324_2 CB@34_mAd325_1 CB@34_mAd325_2 CB@34_mAd326_1 CB@34_mAd326_2 CB@34_mAd327_1 CB@34_mAd327_2 CB@34_mAd330_1 CB@34_mAd330_2 CB@34_mAd331_1 CB@34_mAd331_2 CB@34_mAd332_1 CB@34_mAd332_2 CB@34_mAd333_1 
+CB@34_mAd333_2 CB@34_mAd334_1 CB@34_mAd334_2 CB@34_mAd335_1 CB@34_mAd335_2 CB@34_mAd336_1 CB@34_mAd336_2 CB@34_mAd337_1 CB@34_mAd337_2 CB@34_mAd340_1 CB@34_mAd340_2 CB@34_mAd341_1 CB@34_mAd341_2 CB@34_mAd342_1 CB@34_mAd342_2 CB@34_mAd343_1 CB@34_mAd343_2 CB@34_mAd344_1 CB@34_mAd344_2 CB@34_mAd345_1 CB@34_mAd345_2 CB@34_mAd346_1 CB@34_mAd346_2 CB@34_mAd347_1 CB@34_mAd347_2 CB@34_mAd350_1 CB@34_mAd350_2 CB@34_mAd351_1 CB@34_mAd351_2 CB@34_mAd352_1 CB@34_mAd352_2 CB@34_mAd353_1 CB@34_mAd353_2 CB@34_mAd354_1 
+CB@34_mAd354_2 CB@34_mAd355_1 CB@34_mAd355_2 CB@34_mAd356_1 CB@34_mAd356_2 CB@34_mAd357_1 CB@34_mAd357_2 CB@34_mAd360_1 CB@34_mAd360_2 CB@34_mAd361_1 CB@34_mAd361_2 CB@34_mAd362_1 CB@34_mAd362_2 CB@34_mAd363_1 CB@34_mAd363_2 CB@34_mAd364_1 CB@34_mAd364_2 CB@34_mAd365_1 CB@34_mAd365_2 CB@34_mAd366_1 CB@34_mAd366_2 CB@34_mAd367_1 CB@34_mAd367_2 CB@34_mAd371_1 CB@34_mAd371_2 CB@34_mAd372_1 CB@34_mAd372_2 CB@34_mAd373_1 CB@34_mAd373_2 CB@34_mAd374_1 CB@34_mAd374_2 CB@34_mAd375_1 CB@34_mAd375_2 CB@34_mAd376_1 
+CB@34_mAd376_2 CB@34_mAd377_1 CB@34_mAd377_2 CB@34_mAd400_1 CB@34_mAd400_2 CB@34_mAd401_1 CB@34_mAd401_2 CB@34_mAd402_1 CB@34_mAd402_2 CB@34_mAd403_1 CB@34_mAd403_2 CB@34_mAd404_1 CB@34_mAd404_2 CB@34_mAd405_1 CB@34_mAd405_2 CB@34_mAd406_1 CB@34_mAd406_2 CB@34_mAd407_1 CB@34_mAd407_2 CB@34_mAd410_1 CB@34_mAd410_2 CB@34_mAd411_1 CB@34_mAd411_2 CB@34_mAd412_1 CB@34_mAd412_2 CB@34_mAd413_1 CB@34_mAd413_2 CB@34_mAd414_1 CB@34_mAd414_2 CB@34_mAd415_1 CB@34_mAd415_2 CB@34_mAd416_1 CB@34_mAd416_2 CB@34_mAd417_1 
+CB@34_mAd417_2 CB@34_mAd420_1 CB@34_mAd420_2 CB@34_mAd421_1 CB@34_mAd421_2 CB@34_mAd422_1 CB@34_mAd422_2 CB@34_mAd423_1 CB@34_mAd423_2 CB@34_mAd424_1 CB@34_mAd424_2 CB@34_mAd425_1 CB@34_mAd425_2 CB@34_mAd426_1 CB@34_mAd426_2 CB@34_mAd427_1 CB@34_mAd427_2 CB@34_mAd430_1 CB@34_mAd430_2 CB@34_mAd431_1 CB@34_mAd431_2 CB@34_mAd432_1 CB@34_mAd432_2 CB@34_mAd433_1 CB@34_mAd433_2 CB@34_mAd434_1 CB@34_mAd434_2 CB@34_mAd435_1 CB@34_mAd435_2 CB@34_mAd436_1 CB@34_mAd436_2 CB@34_mAd437_1 CB@34_mAd437_2 CB@34_mAd440_1 
+CB@34_mAd440_2 CB@34_mAd441_1 CB@34_mAd441_2 CB@34_mAd442_1 CB@34_mAd442_2 CB@34_mAd443_1 CB@34_mAd443_2 CB@34_mAd444_1 CB@34_mAd444_2 CB@34_mAd445_1 CB@34_mAd445_2 CB@34_mAd446_1 CB@34_mAd446_2 CB@34_mAd447_1 CB@34_mAd447_2 CB@34_mAd450_1 CB@34_mAd450_2 CB@34_mAd451_1 CB@34_mAd451_2 CB@34_mAd452_1 CB@34_mAd452_2 CB@34_mAd453_1 CB@34_mAd453_2 CB@34_mAd454_1 CB@34_mAd454_2 CB@34_mAd455_1 CB@34_mAd455_2 CB@34_mAd456_1 CB@34_mAd456_2 CB@34_mAd457_1 CB@34_mAd457_2 CB@34_mAd460_1 CB@34_mAd460_2 CB@34_mAd466_1 
+CB@34_mAd466_2 CB@34_mAd467_1 CB@34_mAd467_2 CB@34_mAd500_1 CB@34_mAd500_2 CB@34_mAd501_1 CB@34_mAd501_2 CB@34_mAd502_1 CB@34_mAd502_2 CB@34_mAd508_1 CB@34_mAd508_2 CB@34_mAd509_1 CB@34_mAd509_2 CB@34_mAd512_1 CB@34_mAd512_2 CB@34_mAd513_1 CB@34_mAd513_2 CB@34_mAd514_1 CB@34_mAd514_2 CB@34_mAd515_1 CB@34_mAd515_2 CB@34_mAd516_1 CB@34_mAd516_2 CB@34_mAd517_1 CB@34_mAd517_2 CB@34_mAd520_1 CB@34_mAd520_2 CB@34_mAd521_1 CB@34_mAd521_2 CB@34_mAd522_1 CB@34_mAd522_2 CB@34_mAd523_1 CB@34_mAd523_2 CB@34_mAd524_1 
+CB@34_mAd524_2 CB@34_mAd525_1 CB@34_mAd525_2 CB@34_mAd526_1 CB@34_mAd526_2 CB@34_mAd527_1 CB@34_mAd527_2 CB@34_mAd530_1 CB@34_mAd530_2 CB@34_mAd531_1 CB@34_mAd531_2 CB@34_mAd532_1 CB@34_mAd532_2 CB@34_mAd533_1 CB@34_mAd533_2 CB@34_mAd534_1 CB@34_mAd534_2 CB@34_mAd535_1 CB@34_mAd535_2 CB@34_mAd536_1 CB@34_mAd536_2 CB@34_mAd537_1 CB@34_mAd537_2 CB@34_mAd540_1 CB@34_mAd540_2 CB@34_mAd541_1 CB@34_mAd541_2 CB@34_mAd542_1 CB@34_mAd542_2 CB@34_mAd543_1 CB@34_mAd543_2 CB@34_mAd544_1 CB@34_mAd544_2 CB@34_mAd545_1 
+CB@34_mAd545_2 CB@34_mAd546_1 CB@34_mAd546_2 CB@34_mAd547_1 CB@34_mAd547_2 CB@34_mAd550_1 CB@34_mAd550_2 CB@34_mAd551_1 CB@34_mAd551_2 CB@34_mAd552_1 CB@34_mAd552_2 CB@34_mAd553_1 CB@34_mAd553_2 CB@34_mAd554_1 CB@34_mAd554_2 CB@34_mAd555_1 CB@34_mAd555_2 CB@34_mAd556_1 CB@34_mAd556_2 CB@34_mAd557_1 CB@34_mAd557_2 CB@34_mAd560_1 CB@34_mAd560_2 CB@34_mAd561_1 CB@34_mAd561_2 CB@34_mAd562_1 CB@34_mAd562_2 CB@34_mAd563_1 CB@34_mAd563_2 CB@34_mAd564_1 CB@34_mAd564_2 CB@34_mAd565_1 CB@34_mAd565_2 CB@34_mAd566_1 
+CB@34_mAd566_2 CB@34_mAd567_1 CB@34_mAd567_2 CB@34_mAd570_1 CB@34_mAd570_2 CB@34_mAd571_1 CB@34_mAd571_2 CB@34_mAd572_1 CB@34_mAd572_2 CB@34_mAd573_1 CB@34_mAd573_2 CB@34_mAd575_1 CB@34_mAd575_2 CB@34_mAd576_1 CB@34_mAd576_2 CB@34_mAd577_1 CB@34_mAd577_2 CB@34_mAd600_1 CB@34_mAd600_2 CB@34_mAd601_1 CB@34_mAd601_2 CB@34_mAd602_1 CB@34_mAd602_2 CB@34_mAd604_1 CB@34_mAd604_2 CB@34_mAd605_1 CB@34_mAd605_2 CB@34_mAd606_1 CB@34_mAd606_2 CB@34_mAd607_1 CB@34_mAd607_2 CB@34_mAd610_1 CB@34_mAd610_2 CB@34_mAd611_1 
+CB@34_mAd611_2 CB@34_mAd612_1 CB@34_mAd612_2 CB@34_mAd613_1 CB@34_mAd613_2 CB@34_mAd614_1 CB@34_mAd614_2 CB@34_mAd615_1 CB@34_mAd615_2 CB@34_mAd616_1 CB@34_mAd616_2 CB@34_mAd617_1 CB@34_mAd617_2 CB@34_mAd620_1 CB@34_mAd620_2 CB@34_mAd621_1 CB@34_mAd621_2 CB@34_mAd622_1 CB@34_mAd622_2 CB@34_mAd623_1 CB@34_mAd623_2 CB@34_mAd624_1 CB@34_mAd624_2 CB@34_mAd625_1 CB@34_mAd625_2 CB@34_mAd626_1 CB@34_mAd626_2 CB@34_mAd627_1 CB@34_mAd627_2 CB@34_mAd630_1 CB@34_mAd630_2 CB@34_mAd631_1 CB@34_mAd631_2 CB@34_mAd632_1 
+CB@34_mAd632_2 CB@34_mAd633_1 CB@34_mAd633_2 CB@34_mAd634_1 CB@34_mAd634_2 CB@34_mAd635_1 CB@34_mAd635_2 CB@34_mAd636_1 CB@34_mAd636_2 CB@34_mAd637_1 CB@34_mAd637_2 CB@34_mAd640_1 CB@34_mAd640_2 CB@34_mAd641_1 CB@34_mAd641_2 CB@34_mAd642_1 CB@34_mAd642_2 CB@34_mAd643_1 CB@34_mAd643_2 CB@34_mAd644_1 CB@34_mAd644_2 CB@34_mAd645_1 CB@34_mAd645_2 CB@34_mAd646_1 CB@34_mAd646_2 CB@34_mAd647_1 CB@34_mAd647_2 CB@34_mAd650_1 CB@34_mAd650_2 CB@34_mAd651_1 CB@34_mAd651_2 CB@34_mAd652_1 CB@34_mAd652_2 CB@34_mAd653_1 
+CB@34_mAd653_2 CB@34_mAd654_1 CB@34_mAd654_2 CB@34_mAd655_1 CB@34_mAd655_2 CB@34_mAd656_1 CB@34_mAd656_2 CB@34_mAd657_1 CB@34_mAd657_2 CB@34_mAd660_1 CB@34_mAd660_2 CB@34_mAd661_1 CB@34_mAd661_2 CB@34_mAd662_1 CB@34_mAd662_2 CB@34_mAd663_1 CB@34_mAd663_2 CB@34_mAd664_1 CB@34_mAd664_2 CB@34_mAd665_1 CB@34_mAd665_2 CB@34_mAd666_1 CB@34_mAd666_2 CB@34_mAd667_1 CB@34_mAd667_2 CB@34_mAd675_1 CB@34_mAd675_2 CB@34_mAd676_1 CB@34_mAd676_2 CB@34_mAd677_1 CB@34_mAd677_2 CB@34_mAd700_1 CB@34_mAd700_2 CB@34_mAd710_1 
+CB@34_mAd710_2 CB@34_mAd711_1 CB@34_mAd711_2 CB@34_mAd717_1 CB@34_mAd717_2 CB@34_mAd720_1 CB@34_mAd720_2 CB@34_mAd721_1 CB@34_mAd721_2 CB@34_mAd722_1 CB@34_mAd722_2 CB@34_mAd723_1 CB@34_mAd723_2 CB@34_mAd724_1 CB@34_mAd724_2 CB@34_mAd725_1 CB@34_mAd725_2 CB@34_mAd726_1 CB@34_mAd726_2 CB@34_mAd727_1 CB@34_mAd727_2 CB@34_mAd730_1 CB@34_mAd730_2 CB@34_mAd731_1 CB@34_mAd731_2 CB@34_mAd732_1 CB@34_mAd732_2 CB@34_mAd733_1 CB@34_mAd733_2 CB@34_mAd734_1 CB@34_mAd734_2 CB@34_mAd735_1 CB@34_mAd735_2 CB@34_mAd736_1 
+CB@34_mAd736_2 CB@34_mAd737_1 CB@34_mAd737_2 CB@34_mAd740_1 CB@34_mAd740_2 CB@34_mAd741_1 CB@34_mAd741_2 CB@34_mAd742_1 CB@34_mAd742_2 CB@34_mAd743_1 CB@34_mAd743_2 CB@34_mAd744_1 CB@34_mAd744_2 CB@34_mAd745_1 CB@34_mAd745_2 CB@34_mAd746_1 CB@34_mAd746_2 CB@34_mAd747_1 CB@34_mAd747_2 CB@34_mAd750_1 CB@34_mAd750_2 CB@34_mAd751_1 CB@34_mAd751_2 CB@34_mAd752_1 CB@34_mAd752_2 CB@34_mAd753_1 CB@34_mAd753_2 CB@34_mAd754_1 CB@34_mAd754_2 CB@34_mAd755_1 CB@34_mAd755_2 CB@34_mAd756_1 CB@34_mAd756_2 CB@34_mAd757_1 
+CB@34_mAd757_2 CB@34_mAd760_1 CB@34_mAd760_2 CB@34_mAd761_1 CB@34_mAd761_2 CB@34_mAd762_1 CB@34_mAd762_2 CB@34_mAd763_1 CB@34_mAd763_2 CB@34_mAd764_1 CB@34_mAd764_2 CB@34_mAd765_1 CB@34_mAd765_2 CB@34_mAd766_1 CB@34_mAd766_2 CB@34_mAd767_1 CB@34_mAd767_2 CB@34_mAd771_1 CB@34_mAd771_2 CB@34_mAd772_1 CB@34_mAd772_2 CB@34_mAd773_1 CB@34_mAd773_2 CB@34_mAd774_1 CB@34_mAd774_2 CB@34_mAd775_1 CB@34_mAd775_2 CB@34_mAd776_1 CB@34_mAd776_2 CB@34_mAd777_1 CB@34_mAd777_2 CB@34_X0 CB@34_X1 CB@34_X10 CB@34_X11 
+CB@34_X12 CB@34_X13 CB@34_X2 CB@34_X3 CB@34_X4 CB@34_X5 CB@34_X6 CB@34_X7 CB@34_X8 CB@34_X9 CB@34_Y1 CB@34_Y10 CB@34_Y11 CB@34_Y12 CB@34_Y2 CB@34_Y3 CB@34_Y4 CB@34_Y5 CB@34_Y6 CB@34_Y7 CB@34_Y8 CB@34_Y9 CB@34_Z1 CB@34_Z10 CB@34_Z11 CB@34_Z12 CB@34_Z2 CB@34_Z3 CB@34_Z4 CB@34_Z5 CB@34_Z6 CB@34_Z7 CB@34_Z8 CB@34_Z9 _5400TP094__CB
XCB@35 CB@35_K0 CB@35_K1 CB@35_K10 CB@35_K11 CB@35_K12 CB@35_K13 CB@35_K2 CB@35_K3 CB@35_K4 CB@35_K5 CB@35_K6 CB@35_K7 CB@35_K8 CB@35_K9 CB@35_mAd000_1 CB@35_mAd000_2 CB@35_mAd001_1 CB@35_mAd001_2 CB@35_mAd002_1 CB@35_mAd002_2 CB@35_mAd003_1 CB@35_mAd003_2 CB@35_mAd004_1 CB@35_mAd004_2 CB@35_mAd005_1 CB@35_mAd005_2 CB@35_mAd006_1 CB@35_mAd006_2 CB@35_mAd007_1 CB@35_mAd007_2 CB@35_mAd010_1 CB@35_mAd010_2 CB@35_mAd011_1 CB@35_mAd011_2 CB@35_mAd012_1 CB@35_mAd012_2 CB@35_mAd013_1 CB@35_mAd013_2 CB@35_mAd014_1 
+CB@35_mAd014_2 CB@35_mAd015_1 CB@35_mAd015_2 CB@35_mAd016_1 CB@35_mAd016_2 CB@35_mAd017_1 CB@35_mAd017_2 CB@35_mAd020_1 CB@35_mAd020_2 CB@35_mAd021_1 CB@35_mAd021_2 CB@35_mAd022_1 CB@35_mAd022_2 CB@35_mAd023_1 CB@35_mAd023_2 CB@35_mAd024_1 CB@35_mAd024_2 CB@35_mAd025_1 CB@35_mAd025_2 CB@35_mAd026_1 CB@35_mAd026_2 CB@35_mAd027_1 CB@35_mAd027_2 CB@35_mAd030_1 CB@35_mAd030_2 CB@35_mAd031_1 CB@35_mAd031_2 CB@35_mAd032_1 CB@35_mAd032_2 CB@35_mAd033_1 CB@35_mAd033_2 CB@35_mAd034_1 CB@35_mAd034_2 CB@35_mAd035_1 
+CB@35_mAd035_2 CB@35_mAd036_1 CB@35_mAd036_2 CB@35_mAd037_1 CB@35_mAd037_2 CB@35_mAd040_1 CB@35_mAd040_2 CB@35_mAd041_1 CB@35_mAd041_2 CB@35_mAd042_1 CB@35_mAd042_2 CB@35_mAd043_1 CB@35_mAd043_2 CB@35_mAd044_1 CB@35_mAd044_2 CB@35_mAd045_1 CB@35_mAd045_2 CB@35_mAd046_1 CB@35_mAd046_2 CB@35_mAd047_1 CB@35_mAd047_2 CB@35_mAd050_1 CB@35_mAd050_2 CB@35_mAd051_1 CB@35_mAd051_2 CB@35_mAd052_1 CB@35_mAd052_2 CB@35_mAd053_1 CB@35_mAd053_2 CB@35_mAd054_1 CB@35_mAd054_2 CB@35_mAd055_1 CB@35_mAd055_2 CB@35_mAd056_1 
+CB@35_mAd056_2 CB@35_mAd057_1 CB@35_mAd057_2 CB@35_mAd060_1 CB@35_mAd060_2 CB@35_mAd066_1 CB@35_mAd066_2 CB@35_mAd067_1 CB@35_mAd067_2 CB@35_mAd100_1 CB@35_mAd100_2 CB@35_mAd101_1 CB@35_mAd101_2 CB@35_mAd102_1 CB@35_mAd102_2 CB@35_mAd110_1 CB@35_mAd110_2 CB@35_mAd111_1 CB@35_mAd111_2 CB@35_mAd112_1 CB@35_mAd112_2 CB@35_mAd113_1 CB@35_mAd113_2 CB@35_mAd114_1 CB@35_mAd114_2 CB@35_mAd115_1 CB@35_mAd115_2 CB@35_mAd116_1 CB@35_mAd116_2 CB@35_mAd117_1 CB@35_mAd117_2 CB@35_mAd120_1 CB@35_mAd120_2 CB@35_mAd121_1 
+CB@35_mAd121_2 CB@35_mAd122_1 CB@35_mAd122_2 CB@35_mAd123_1 CB@35_mAd123_2 CB@35_mAd124_1 CB@35_mAd124_2 CB@35_mAd125_1 CB@35_mAd125_2 CB@35_mAd126_1 CB@35_mAd126_2 CB@35_mAd127_1 CB@35_mAd127_2 CB@35_mAd130_1 CB@35_mAd130_2 CB@35_mAd131_1 CB@35_mAd131_2 CB@35_mAd132_1 CB@35_mAd132_2 CB@35_mAd133_1 CB@35_mAd133_2 CB@35_mAd134_1 CB@35_mAd134_2 CB@35_mAd135_1 CB@35_mAd135_2 CB@35_mAd136_1 CB@35_mAd136_2 CB@35_mAd137_1 CB@35_mAd137_2 CB@35_mAd140_1 CB@35_mAd140_2 CB@35_mAd141_1 CB@35_mAd141_2 CB@35_mAd142_1 
+CB@35_mAd142_2 CB@35_mAd143_1 CB@35_mAd143_2 CB@35_mAd144_1 CB@35_mAd144_2 CB@35_mAd145_1 CB@35_mAd145_2 CB@35_mAd146_1 CB@35_mAd146_2 CB@35_mAd147_1 CB@35_mAd147_2 CB@35_mAd150_1 CB@35_mAd150_2 CB@35_mAd151_1 CB@35_mAd151_2 CB@35_mAd152_1 CB@35_mAd152_2 CB@35_mAd153_1 CB@35_mAd153_2 CB@35_mAd154_1 CB@35_mAd154_2 CB@35_mAd155_1 CB@35_mAd155_2 CB@35_mAd156_1 CB@35_mAd156_2 CB@35_mAd157_1 CB@35_mAd157_2 CB@35_mAd160_1 CB@35_mAd160_2 CB@35_mAd161_1 CB@35_mAd161_2 CB@35_mAd162_1 CB@35_mAd162_2 CB@35_mAd163_1 
+CB@35_mAd163_2 CB@35_mAd164_1 CB@35_mAd164_2 CB@35_mAd165_1 CB@35_mAd165_2 CB@35_mAd166_1 CB@35_mAd166_2 CB@35_mAd167_1 CB@35_mAd167_2 CB@35_mAd170_1 CB@35_mAd170_2 CB@35_mAd171_1 CB@35_mAd171_2 CB@35_mAd172_1 CB@35_mAd172_2 CB@35_mAd173_1 CB@35_mAd173_2 CB@35_mAd175_1 CB@35_mAd175_2 CB@35_mAd176_1 CB@35_mAd176_2 CB@35_mAd177_1 CB@35_mAd177_2 CB@35_mAd200_1 CB@35_mAd200_2 CB@35_mAd201_1 CB@35_mAd201_2 CB@35_mAd202_1 CB@35_mAd202_2 CB@35_mAd204_1 CB@35_mAd204_2 CB@35_mAd205_1 CB@35_mAd205_2 CB@35_mAd206_1 
+CB@35_mAd206_2 CB@35_mAd207_1 CB@35_mAd207_2 CB@35_mAd210_1 CB@35_mAd210_2 CB@35_mAd211_1 CB@35_mAd211_2 CB@35_mAd212_1 CB@35_mAd212_2 CB@35_mAd213_1 CB@35_mAd213_2 CB@35_mAd214_1 CB@35_mAd214_2 CB@35_mAd215_1 CB@35_mAd215_2 CB@35_mAd216_1 CB@35_mAd216_2 CB@35_mAd217_1 CB@35_mAd217_2 CB@35_mAd220_1 CB@35_mAd220_2 CB@35_mAd221_1 CB@35_mAd221_2 CB@35_mAd222_1 CB@35_mAd222_2 CB@35_mAd223_1 CB@35_mAd223_2 CB@35_mAd224_1 CB@35_mAd224_2 CB@35_mAd225_1 CB@35_mAd225_2 CB@35_mAd226_1 CB@35_mAd226_2 CB@35_mAd227_1 
+CB@35_mAd227_2 CB@35_mAd230_1 CB@35_mAd230_2 CB@35_mAd231_1 CB@35_mAd231_2 CB@35_mAd232_1 CB@35_mAd232_2 CB@35_mAd233_1 CB@35_mAd233_2 CB@35_mAd234_1 CB@35_mAd234_2 CB@35_mAd235_1 CB@35_mAd235_2 CB@35_mAd236_1 CB@35_mAd236_2 CB@35_mAd237_1 CB@35_mAd237_2 CB@35_mAd240_1 CB@35_mAd240_2 CB@35_mAd241_1 CB@35_mAd241_2 CB@35_mAd242_1 CB@35_mAd242_2 CB@35_mAd243_1 CB@35_mAd243_2 CB@35_mAd244_1 CB@35_mAd244_2 CB@35_mAd245_1 CB@35_mAd245_2 CB@35_mAd246_1 CB@35_mAd246_2 CB@35_mAd247_1 CB@35_mAd247_2 CB@35_mAd250_1 
+CB@35_mAd250_2 CB@35_mAd251_1 CB@35_mAd251_2 CB@35_mAd252_1 CB@35_mAd252_2 CB@35_mAd253_1 CB@35_mAd253_2 CB@35_mAd254_1 CB@35_mAd254_2 CB@35_mAd255_1 CB@35_mAd255_2 CB@35_mAd256_1 CB@35_mAd256_2 CB@35_mAd257_1 CB@35_mAd257_2 CB@35_mAd260_1 CB@35_mAd260_2 CB@35_mAd261_1 CB@35_mAd261_2 CB@35_mAd262_1 CB@35_mAd262_2 CB@35_mAd263_1 CB@35_mAd263_2 CB@35_mAd264_1 CB@35_mAd264_2 CB@35_mAd265_1 CB@35_mAd265_2 CB@35_mAd266_1 CB@35_mAd266_2 CB@35_mAd267_1 CB@35_mAd267_2 CB@35_mAd275_1 CB@35_mAd275_2 CB@35_mAd276_1 
+CB@35_mAd276_2 CB@35_mAd277_1 CB@35_mAd277_2 CB@35_mAd300_1 CB@35_mAd300_2 CB@35_mAd310_1 CB@35_mAd310_2 CB@35_mAd311_1 CB@35_mAd311_2 CB@35_mAd317_1 CB@35_mAd317_2 CB@35_mAd320_1 CB@35_mAd320_2 CB@35_mAd321_1 CB@35_mAd321_2 CB@35_mAd322_1 CB@35_mAd322_2 CB@35_mAd323_1 CB@35_mAd323_2 CB@35_mAd324_1 CB@35_mAd324_2 CB@35_mAd325_1 CB@35_mAd325_2 CB@35_mAd326_1 CB@35_mAd326_2 CB@35_mAd327_1 CB@35_mAd327_2 CB@35_mAd330_1 CB@35_mAd330_2 CB@35_mAd331_1 CB@35_mAd331_2 CB@35_mAd332_1 CB@35_mAd332_2 CB@35_mAd333_1 
+CB@35_mAd333_2 CB@35_mAd334_1 CB@35_mAd334_2 CB@35_mAd335_1 CB@35_mAd335_2 CB@35_mAd336_1 CB@35_mAd336_2 CB@35_mAd337_1 CB@35_mAd337_2 CB@35_mAd340_1 CB@35_mAd340_2 CB@35_mAd341_1 CB@35_mAd341_2 CB@35_mAd342_1 CB@35_mAd342_2 CB@35_mAd343_1 CB@35_mAd343_2 CB@35_mAd344_1 CB@35_mAd344_2 CB@35_mAd345_1 CB@35_mAd345_2 CB@35_mAd346_1 CB@35_mAd346_2 CB@35_mAd347_1 CB@35_mAd347_2 CB@35_mAd350_1 CB@35_mAd350_2 CB@35_mAd351_1 CB@35_mAd351_2 CB@35_mAd352_1 CB@35_mAd352_2 CB@35_mAd353_1 CB@35_mAd353_2 CB@35_mAd354_1 
+CB@35_mAd354_2 CB@35_mAd355_1 CB@35_mAd355_2 CB@35_mAd356_1 CB@35_mAd356_2 CB@35_mAd357_1 CB@35_mAd357_2 CB@35_mAd360_1 CB@35_mAd360_2 CB@35_mAd361_1 CB@35_mAd361_2 CB@35_mAd362_1 CB@35_mAd362_2 CB@35_mAd363_1 CB@35_mAd363_2 CB@35_mAd364_1 CB@35_mAd364_2 CB@35_mAd365_1 CB@35_mAd365_2 CB@35_mAd366_1 CB@35_mAd366_2 CB@35_mAd367_1 CB@35_mAd367_2 CB@35_mAd371_1 CB@35_mAd371_2 CB@35_mAd372_1 CB@35_mAd372_2 CB@35_mAd373_1 CB@35_mAd373_2 CB@35_mAd374_1 CB@35_mAd374_2 CB@35_mAd375_1 CB@35_mAd375_2 CB@35_mAd376_1 
+CB@35_mAd376_2 CB@35_mAd377_1 CB@35_mAd377_2 CB@35_mAd400_1 CB@35_mAd400_2 CB@35_mAd401_1 CB@35_mAd401_2 CB@35_mAd402_1 CB@35_mAd402_2 CB@35_mAd403_1 CB@35_mAd403_2 CB@35_mAd404_1 CB@35_mAd404_2 CB@35_mAd405_1 CB@35_mAd405_2 CB@35_mAd406_1 CB@35_mAd406_2 CB@35_mAd407_1 CB@35_mAd407_2 CB@35_mAd410_1 CB@35_mAd410_2 CB@35_mAd411_1 CB@35_mAd411_2 CB@35_mAd412_1 CB@35_mAd412_2 CB@35_mAd413_1 CB@35_mAd413_2 CB@35_mAd414_1 CB@35_mAd414_2 CB@35_mAd415_1 CB@35_mAd415_2 CB@35_mAd416_1 CB@35_mAd416_2 CB@35_mAd417_1 
+CB@35_mAd417_2 CB@35_mAd420_1 CB@35_mAd420_2 CB@35_mAd421_1 CB@35_mAd421_2 CB@35_mAd422_1 CB@35_mAd422_2 CB@35_mAd423_1 CB@35_mAd423_2 CB@35_mAd424_1 CB@35_mAd424_2 CB@35_mAd425_1 CB@35_mAd425_2 CB@35_mAd426_1 CB@35_mAd426_2 CB@35_mAd427_1 CB@35_mAd427_2 CB@35_mAd430_1 CB@35_mAd430_2 CB@35_mAd431_1 CB@35_mAd431_2 CB@35_mAd432_1 CB@35_mAd432_2 CB@35_mAd433_1 CB@35_mAd433_2 CB@35_mAd434_1 CB@35_mAd434_2 CB@35_mAd435_1 CB@35_mAd435_2 CB@35_mAd436_1 CB@35_mAd436_2 CB@35_mAd437_1 CB@35_mAd437_2 CB@35_mAd440_1 
+CB@35_mAd440_2 CB@35_mAd441_1 CB@35_mAd441_2 CB@35_mAd442_1 CB@35_mAd442_2 CB@35_mAd443_1 CB@35_mAd443_2 CB@35_mAd444_1 CB@35_mAd444_2 CB@35_mAd445_1 CB@35_mAd445_2 CB@35_mAd446_1 CB@35_mAd446_2 CB@35_mAd447_1 CB@35_mAd447_2 CB@35_mAd450_1 CB@35_mAd450_2 CB@35_mAd451_1 CB@35_mAd451_2 CB@35_mAd452_1 CB@35_mAd452_2 CB@35_mAd453_1 CB@35_mAd453_2 CB@35_mAd454_1 CB@35_mAd454_2 CB@35_mAd455_1 CB@35_mAd455_2 CB@35_mAd456_1 CB@35_mAd456_2 CB@35_mAd457_1 CB@35_mAd457_2 CB@35_mAd460_1 CB@35_mAd460_2 CB@35_mAd466_1 
+CB@35_mAd466_2 CB@35_mAd467_1 CB@35_mAd467_2 CB@35_mAd500_1 CB@35_mAd500_2 CB@35_mAd501_1 CB@35_mAd501_2 CB@35_mAd502_1 CB@35_mAd502_2 CB@35_mAd508_1 CB@35_mAd508_2 CB@35_mAd509_1 CB@35_mAd509_2 CB@35_mAd512_1 CB@35_mAd512_2 CB@35_mAd513_1 CB@35_mAd513_2 CB@35_mAd514_1 CB@35_mAd514_2 CB@35_mAd515_1 CB@35_mAd515_2 CB@35_mAd516_1 CB@35_mAd516_2 CB@35_mAd517_1 CB@35_mAd517_2 CB@35_mAd520_1 CB@35_mAd520_2 CB@35_mAd521_1 CB@35_mAd521_2 CB@35_mAd522_1 CB@35_mAd522_2 CB@35_mAd523_1 CB@35_mAd523_2 CB@35_mAd524_1 
+CB@35_mAd524_2 CB@35_mAd525_1 CB@35_mAd525_2 CB@35_mAd526_1 CB@35_mAd526_2 CB@35_mAd527_1 CB@35_mAd527_2 CB@35_mAd530_1 CB@35_mAd530_2 CB@35_mAd531_1 CB@35_mAd531_2 CB@35_mAd532_1 CB@35_mAd532_2 CB@35_mAd533_1 CB@35_mAd533_2 CB@35_mAd534_1 CB@35_mAd534_2 CB@35_mAd535_1 CB@35_mAd535_2 CB@35_mAd536_1 CB@35_mAd536_2 CB@35_mAd537_1 CB@35_mAd537_2 CB@35_mAd540_1 CB@35_mAd540_2 CB@35_mAd541_1 CB@35_mAd541_2 CB@35_mAd542_1 CB@35_mAd542_2 CB@35_mAd543_1 CB@35_mAd543_2 CB@35_mAd544_1 CB@35_mAd544_2 CB@35_mAd545_1 
+CB@35_mAd545_2 CB@35_mAd546_1 CB@35_mAd546_2 CB@35_mAd547_1 CB@35_mAd547_2 CB@35_mAd550_1 CB@35_mAd550_2 CB@35_mAd551_1 CB@35_mAd551_2 CB@35_mAd552_1 CB@35_mAd552_2 CB@35_mAd553_1 CB@35_mAd553_2 CB@35_mAd554_1 CB@35_mAd554_2 CB@35_mAd555_1 CB@35_mAd555_2 CB@35_mAd556_1 CB@35_mAd556_2 CB@35_mAd557_1 CB@35_mAd557_2 CB@35_mAd560_1 CB@35_mAd560_2 CB@35_mAd561_1 CB@35_mAd561_2 CB@35_mAd562_1 CB@35_mAd562_2 CB@35_mAd563_1 CB@35_mAd563_2 CB@35_mAd564_1 CB@35_mAd564_2 CB@35_mAd565_1 CB@35_mAd565_2 CB@35_mAd566_1 
+CB@35_mAd566_2 CB@35_mAd567_1 CB@35_mAd567_2 CB@35_mAd570_1 CB@35_mAd570_2 CB@35_mAd571_1 CB@35_mAd571_2 CB@35_mAd572_1 CB@35_mAd572_2 CB@35_mAd573_1 CB@35_mAd573_2 CB@35_mAd575_1 CB@35_mAd575_2 CB@35_mAd576_1 CB@35_mAd576_2 CB@35_mAd577_1 CB@35_mAd577_2 CB@35_mAd600_1 CB@35_mAd600_2 CB@35_mAd601_1 CB@35_mAd601_2 CB@35_mAd602_1 CB@35_mAd602_2 CB@35_mAd604_1 CB@35_mAd604_2 CB@35_mAd605_1 CB@35_mAd605_2 CB@35_mAd606_1 CB@35_mAd606_2 CB@35_mAd607_1 CB@35_mAd607_2 CB@35_mAd610_1 CB@35_mAd610_2 CB@35_mAd611_1 
+CB@35_mAd611_2 CB@35_mAd612_1 CB@35_mAd612_2 CB@35_mAd613_1 CB@35_mAd613_2 CB@35_mAd614_1 CB@35_mAd614_2 CB@35_mAd615_1 CB@35_mAd615_2 CB@35_mAd616_1 CB@35_mAd616_2 CB@35_mAd617_1 CB@35_mAd617_2 CB@35_mAd620_1 CB@35_mAd620_2 CB@35_mAd621_1 CB@35_mAd621_2 CB@35_mAd622_1 CB@35_mAd622_2 CB@35_mAd623_1 CB@35_mAd623_2 CB@35_mAd624_1 CB@35_mAd624_2 CB@35_mAd625_1 CB@35_mAd625_2 CB@35_mAd626_1 CB@35_mAd626_2 CB@35_mAd627_1 CB@35_mAd627_2 CB@35_mAd630_1 CB@35_mAd630_2 CB@35_mAd631_1 CB@35_mAd631_2 CB@35_mAd632_1 
+CB@35_mAd632_2 CB@35_mAd633_1 CB@35_mAd633_2 CB@35_mAd634_1 CB@35_mAd634_2 CB@35_mAd635_1 CB@35_mAd635_2 CB@35_mAd636_1 CB@35_mAd636_2 CB@35_mAd637_1 CB@35_mAd637_2 CB@35_mAd640_1 CB@35_mAd640_2 CB@35_mAd641_1 CB@35_mAd641_2 CB@35_mAd642_1 CB@35_mAd642_2 CB@35_mAd643_1 CB@35_mAd643_2 CB@35_mAd644_1 CB@35_mAd644_2 CB@35_mAd645_1 CB@35_mAd645_2 CB@35_mAd646_1 CB@35_mAd646_2 CB@35_mAd647_1 CB@35_mAd647_2 CB@35_mAd650_1 CB@35_mAd650_2 CB@35_mAd651_1 CB@35_mAd651_2 CB@35_mAd652_1 CB@35_mAd652_2 CB@35_mAd653_1 
+CB@35_mAd653_2 CB@35_mAd654_1 CB@35_mAd654_2 CB@35_mAd655_1 CB@35_mAd655_2 CB@35_mAd656_1 CB@35_mAd656_2 CB@35_mAd657_1 CB@35_mAd657_2 CB@35_mAd660_1 CB@35_mAd660_2 CB@35_mAd661_1 CB@35_mAd661_2 CB@35_mAd662_1 CB@35_mAd662_2 CB@35_mAd663_1 CB@35_mAd663_2 CB@35_mAd664_1 CB@35_mAd664_2 CB@35_mAd665_1 CB@35_mAd665_2 CB@35_mAd666_1 CB@35_mAd666_2 CB@35_mAd667_1 CB@35_mAd667_2 CB@35_mAd675_1 CB@35_mAd675_2 CB@35_mAd676_1 CB@35_mAd676_2 CB@35_mAd677_1 CB@35_mAd677_2 CB@35_mAd700_1 CB@35_mAd700_2 CB@35_mAd710_1 
+CB@35_mAd710_2 CB@35_mAd711_1 CB@35_mAd711_2 CB@35_mAd717_1 CB@35_mAd717_2 CB@35_mAd720_1 CB@35_mAd720_2 CB@35_mAd721_1 CB@35_mAd721_2 CB@35_mAd722_1 CB@35_mAd722_2 CB@35_mAd723_1 CB@35_mAd723_2 CB@35_mAd724_1 CB@35_mAd724_2 CB@35_mAd725_1 CB@35_mAd725_2 CB@35_mAd726_1 CB@35_mAd726_2 CB@35_mAd727_1 CB@35_mAd727_2 CB@35_mAd730_1 CB@35_mAd730_2 CB@35_mAd731_1 CB@35_mAd731_2 CB@35_mAd732_1 CB@35_mAd732_2 CB@35_mAd733_1 CB@35_mAd733_2 CB@35_mAd734_1 CB@35_mAd734_2 CB@35_mAd735_1 CB@35_mAd735_2 CB@35_mAd736_1 
+CB@35_mAd736_2 CB@35_mAd737_1 CB@35_mAd737_2 CB@35_mAd740_1 CB@35_mAd740_2 CB@35_mAd741_1 CB@35_mAd741_2 CB@35_mAd742_1 CB@35_mAd742_2 CB@35_mAd743_1 CB@35_mAd743_2 CB@35_mAd744_1 CB@35_mAd744_2 CB@35_mAd745_1 CB@35_mAd745_2 CB@35_mAd746_1 CB@35_mAd746_2 CB@35_mAd747_1 CB@35_mAd747_2 CB@35_mAd750_1 CB@35_mAd750_2 CB@35_mAd751_1 CB@35_mAd751_2 CB@35_mAd752_1 CB@35_mAd752_2 CB@35_mAd753_1 CB@35_mAd753_2 CB@35_mAd754_1 CB@35_mAd754_2 CB@35_mAd755_1 CB@35_mAd755_2 CB@35_mAd756_1 CB@35_mAd756_2 CB@35_mAd757_1 
+CB@35_mAd757_2 CB@35_mAd760_1 CB@35_mAd760_2 CB@35_mAd761_1 CB@35_mAd761_2 CB@35_mAd762_1 CB@35_mAd762_2 CB@35_mAd763_1 CB@35_mAd763_2 CB@35_mAd764_1 CB@35_mAd764_2 CB@35_mAd765_1 CB@35_mAd765_2 CB@35_mAd766_1 CB@35_mAd766_2 CB@35_mAd767_1 CB@35_mAd767_2 CB@35_mAd771_1 CB@35_mAd771_2 CB@35_mAd772_1 CB@35_mAd772_2 CB@35_mAd773_1 CB@35_mAd773_2 CB@35_mAd774_1 CB@35_mAd774_2 CB@35_mAd775_1 CB@35_mAd775_2 CB@35_mAd776_1 CB@35_mAd776_2 CB@35_mAd777_1 CB@35_mAd777_2 CB@35_X0 CB@35_X1 CB@35_X10 CB@35_X11 
+CB@35_X12 CB@35_X13 CB@35_X2 CB@35_X3 CB@35_X4 CB@35_X5 CB@35_X6 CB@35_X7 CB@35_X8 CB@35_X9 CB@35_Y1 CB@35_Y10 CB@35_Y11 CB@35_Y12 CB@35_Y2 CB@35_Y3 CB@35_Y4 CB@35_Y5 CB@35_Y6 CB@35_Y7 CB@35_Y8 CB@35_Y9 CB@35_Z1 CB@35_Z10 CB@35_Z11 CB@35_Z12 CB@35_Z2 CB@35_Z3 CB@35_Z4 CB@35_Z5 CB@35_Z6 CB@35_Z7 CB@35_Z8 CB@35_Z9 _5400TP094__CB
XCB@36 CB@36_K0 CB@36_K1 CB@36_K10 CB@36_K11 CB@36_K12 CB@36_K13 CB@36_K2 CB@36_K3 CB@36_K4 CB@36_K5 CB@36_K6 CB@36_K7 CB@36_K8 CB@36_K9 CB@36_mAd000_1 CB@36_mAd000_2 CB@36_mAd001_1 CB@36_mAd001_2 CB@36_mAd002_1 CB@36_mAd002_2 CB@36_mAd003_1 CB@36_mAd003_2 CB@36_mAd004_1 CB@36_mAd004_2 CB@36_mAd005_1 CB@36_mAd005_2 CB@36_mAd006_1 CB@36_mAd006_2 CB@36_mAd007_1 CB@36_mAd007_2 CB@36_mAd010_1 CB@36_mAd010_2 CB@36_mAd011_1 CB@36_mAd011_2 CB@36_mAd012_1 CB@36_mAd012_2 CB@36_mAd013_1 CB@36_mAd013_2 CB@36_mAd014_1 
+CB@36_mAd014_2 CB@36_mAd015_1 CB@36_mAd015_2 CB@36_mAd016_1 CB@36_mAd016_2 CB@36_mAd017_1 CB@36_mAd017_2 CB@36_mAd020_1 CB@36_mAd020_2 CB@36_mAd021_1 CB@36_mAd021_2 CB@36_mAd022_1 CB@36_mAd022_2 CB@36_mAd023_1 CB@36_mAd023_2 CB@36_mAd024_1 CB@36_mAd024_2 CB@36_mAd025_1 CB@36_mAd025_2 CB@36_mAd026_1 CB@36_mAd026_2 CB@36_mAd027_1 CB@36_mAd027_2 CB@36_mAd030_1 CB@36_mAd030_2 CB@36_mAd031_1 CB@36_mAd031_2 CB@36_mAd032_1 CB@36_mAd032_2 CB@36_mAd033_1 CB@36_mAd033_2 CB@36_mAd034_1 CB@36_mAd034_2 CB@36_mAd035_1 
+CB@36_mAd035_2 CB@36_mAd036_1 CB@36_mAd036_2 CB@36_mAd037_1 CB@36_mAd037_2 CB@36_mAd040_1 CB@36_mAd040_2 CB@36_mAd041_1 CB@36_mAd041_2 CB@36_mAd042_1 CB@36_mAd042_2 CB@36_mAd043_1 CB@36_mAd043_2 CB@36_mAd044_1 CB@36_mAd044_2 CB@36_mAd045_1 CB@36_mAd045_2 CB@36_mAd046_1 CB@36_mAd046_2 CB@36_mAd047_1 CB@36_mAd047_2 CB@36_mAd050_1 CB@36_mAd050_2 CB@36_mAd051_1 CB@36_mAd051_2 CB@36_mAd052_1 CB@36_mAd052_2 CB@36_mAd053_1 CB@36_mAd053_2 CB@36_mAd054_1 CB@36_mAd054_2 CB@36_mAd055_1 CB@36_mAd055_2 CB@36_mAd056_1 
+CB@36_mAd056_2 CB@36_mAd057_1 CB@36_mAd057_2 CB@36_mAd060_1 CB@36_mAd060_2 CB@36_mAd066_1 CB@36_mAd066_2 CB@36_mAd067_1 CB@36_mAd067_2 CB@36_mAd100_1 CB@36_mAd100_2 CB@36_mAd101_1 CB@36_mAd101_2 CB@36_mAd102_1 CB@36_mAd102_2 CB@36_mAd110_1 CB@36_mAd110_2 CB@36_mAd111_1 CB@36_mAd111_2 CB@36_mAd112_1 CB@36_mAd112_2 CB@36_mAd113_1 CB@36_mAd113_2 CB@36_mAd114_1 CB@36_mAd114_2 CB@36_mAd115_1 CB@36_mAd115_2 CB@36_mAd116_1 CB@36_mAd116_2 CB@36_mAd117_1 CB@36_mAd117_2 CB@36_mAd120_1 CB@36_mAd120_2 CB@36_mAd121_1 
+CB@36_mAd121_2 CB@36_mAd122_1 CB@36_mAd122_2 CB@36_mAd123_1 CB@36_mAd123_2 CB@36_mAd124_1 CB@36_mAd124_2 CB@36_mAd125_1 CB@36_mAd125_2 CB@36_mAd126_1 CB@36_mAd126_2 CB@36_mAd127_1 CB@36_mAd127_2 CB@36_mAd130_1 CB@36_mAd130_2 CB@36_mAd131_1 CB@36_mAd131_2 CB@36_mAd132_1 CB@36_mAd132_2 CB@36_mAd133_1 CB@36_mAd133_2 CB@36_mAd134_1 CB@36_mAd134_2 CB@36_mAd135_1 CB@36_mAd135_2 CB@36_mAd136_1 CB@36_mAd136_2 CB@36_mAd137_1 CB@36_mAd137_2 CB@36_mAd140_1 CB@36_mAd140_2 CB@36_mAd141_1 CB@36_mAd141_2 CB@36_mAd142_1 
+CB@36_mAd142_2 CB@36_mAd143_1 CB@36_mAd143_2 CB@36_mAd144_1 CB@36_mAd144_2 CB@36_mAd145_1 CB@36_mAd145_2 CB@36_mAd146_1 CB@36_mAd146_2 CB@36_mAd147_1 CB@36_mAd147_2 CB@36_mAd150_1 CB@36_mAd150_2 CB@36_mAd151_1 CB@36_mAd151_2 CB@36_mAd152_1 CB@36_mAd152_2 CB@36_mAd153_1 CB@36_mAd153_2 CB@36_mAd154_1 CB@36_mAd154_2 CB@36_mAd155_1 CB@36_mAd155_2 CB@36_mAd156_1 CB@36_mAd156_2 CB@36_mAd157_1 CB@36_mAd157_2 CB@36_mAd160_1 CB@36_mAd160_2 CB@36_mAd161_1 CB@36_mAd161_2 CB@36_mAd162_1 CB@36_mAd162_2 CB@36_mAd163_1 
+CB@36_mAd163_2 CB@36_mAd164_1 CB@36_mAd164_2 CB@36_mAd165_1 CB@36_mAd165_2 CB@36_mAd166_1 CB@36_mAd166_2 CB@36_mAd167_1 CB@36_mAd167_2 CB@36_mAd170_1 CB@36_mAd170_2 CB@36_mAd171_1 CB@36_mAd171_2 CB@36_mAd172_1 CB@36_mAd172_2 CB@36_mAd173_1 CB@36_mAd173_2 CB@36_mAd175_1 CB@36_mAd175_2 CB@36_mAd176_1 CB@36_mAd176_2 CB@36_mAd177_1 CB@36_mAd177_2 CB@36_mAd200_1 CB@36_mAd200_2 CB@36_mAd201_1 CB@36_mAd201_2 CB@36_mAd202_1 CB@36_mAd202_2 CB@36_mAd204_1 CB@36_mAd204_2 CB@36_mAd205_1 CB@36_mAd205_2 CB@36_mAd206_1 
+CB@36_mAd206_2 CB@36_mAd207_1 CB@36_mAd207_2 CB@36_mAd210_1 CB@36_mAd210_2 CB@36_mAd211_1 CB@36_mAd211_2 CB@36_mAd212_1 CB@36_mAd212_2 CB@36_mAd213_1 CB@36_mAd213_2 CB@36_mAd214_1 CB@36_mAd214_2 CB@36_mAd215_1 CB@36_mAd215_2 CB@36_mAd216_1 CB@36_mAd216_2 CB@36_mAd217_1 CB@36_mAd217_2 CB@36_mAd220_1 CB@36_mAd220_2 CB@36_mAd221_1 CB@36_mAd221_2 CB@36_mAd222_1 CB@36_mAd222_2 CB@36_mAd223_1 CB@36_mAd223_2 CB@36_mAd224_1 CB@36_mAd224_2 CB@36_mAd225_1 CB@36_mAd225_2 CB@36_mAd226_1 CB@36_mAd226_2 CB@36_mAd227_1 
+CB@36_mAd227_2 CB@36_mAd230_1 CB@36_mAd230_2 CB@36_mAd231_1 CB@36_mAd231_2 CB@36_mAd232_1 CB@36_mAd232_2 CB@36_mAd233_1 CB@36_mAd233_2 CB@36_mAd234_1 CB@36_mAd234_2 CB@36_mAd235_1 CB@36_mAd235_2 CB@36_mAd236_1 CB@36_mAd236_2 CB@36_mAd237_1 CB@36_mAd237_2 CB@36_mAd240_1 CB@36_mAd240_2 CB@36_mAd241_1 CB@36_mAd241_2 CB@36_mAd242_1 CB@36_mAd242_2 CB@36_mAd243_1 CB@36_mAd243_2 CB@36_mAd244_1 CB@36_mAd244_2 CB@36_mAd245_1 CB@36_mAd245_2 CB@36_mAd246_1 CB@36_mAd246_2 CB@36_mAd247_1 CB@36_mAd247_2 CB@36_mAd250_1 
+CB@36_mAd250_2 CB@36_mAd251_1 CB@36_mAd251_2 CB@36_mAd252_1 CB@36_mAd252_2 CB@36_mAd253_1 CB@36_mAd253_2 CB@36_mAd254_1 CB@36_mAd254_2 CB@36_mAd255_1 CB@36_mAd255_2 CB@36_mAd256_1 CB@36_mAd256_2 CB@36_mAd257_1 CB@36_mAd257_2 CB@36_mAd260_1 CB@36_mAd260_2 CB@36_mAd261_1 CB@36_mAd261_2 CB@36_mAd262_1 CB@36_mAd262_2 CB@36_mAd263_1 CB@36_mAd263_2 CB@36_mAd264_1 CB@36_mAd264_2 CB@36_mAd265_1 CB@36_mAd265_2 CB@36_mAd266_1 CB@36_mAd266_2 CB@36_mAd267_1 CB@36_mAd267_2 CB@36_mAd275_1 CB@36_mAd275_2 CB@36_mAd276_1 
+CB@36_mAd276_2 CB@36_mAd277_1 CB@36_mAd277_2 CB@36_mAd300_1 CB@36_mAd300_2 CB@36_mAd310_1 CB@36_mAd310_2 CB@36_mAd311_1 CB@36_mAd311_2 CB@36_mAd317_1 CB@36_mAd317_2 CB@36_mAd320_1 CB@36_mAd320_2 CB@36_mAd321_1 CB@36_mAd321_2 CB@36_mAd322_1 CB@36_mAd322_2 CB@36_mAd323_1 CB@36_mAd323_2 CB@36_mAd324_1 CB@36_mAd324_2 CB@36_mAd325_1 CB@36_mAd325_2 CB@36_mAd326_1 CB@36_mAd326_2 CB@36_mAd327_1 CB@36_mAd327_2 CB@36_mAd330_1 CB@36_mAd330_2 CB@36_mAd331_1 CB@36_mAd331_2 CB@36_mAd332_1 CB@36_mAd332_2 CB@36_mAd333_1 
+CB@36_mAd333_2 CB@36_mAd334_1 CB@36_mAd334_2 CB@36_mAd335_1 CB@36_mAd335_2 CB@36_mAd336_1 CB@36_mAd336_2 CB@36_mAd337_1 CB@36_mAd337_2 CB@36_mAd340_1 CB@36_mAd340_2 CB@36_mAd341_1 CB@36_mAd341_2 CB@36_mAd342_1 CB@36_mAd342_2 CB@36_mAd343_1 CB@36_mAd343_2 CB@36_mAd344_1 CB@36_mAd344_2 CB@36_mAd345_1 CB@36_mAd345_2 CB@36_mAd346_1 CB@36_mAd346_2 CB@36_mAd347_1 CB@36_mAd347_2 CB@36_mAd350_1 CB@36_mAd350_2 CB@36_mAd351_1 CB@36_mAd351_2 CB@36_mAd352_1 CB@36_mAd352_2 CB@36_mAd353_1 CB@36_mAd353_2 CB@36_mAd354_1 
+CB@36_mAd354_2 CB@36_mAd355_1 CB@36_mAd355_2 CB@36_mAd356_1 CB@36_mAd356_2 CB@36_mAd357_1 CB@36_mAd357_2 CB@36_mAd360_1 CB@36_mAd360_2 CB@36_mAd361_1 CB@36_mAd361_2 CB@36_mAd362_1 CB@36_mAd362_2 CB@36_mAd363_1 CB@36_mAd363_2 CB@36_mAd364_1 CB@36_mAd364_2 CB@36_mAd365_1 CB@36_mAd365_2 CB@36_mAd366_1 CB@36_mAd366_2 CB@36_mAd367_1 CB@36_mAd367_2 CB@36_mAd371_1 CB@36_mAd371_2 CB@36_mAd372_1 CB@36_mAd372_2 CB@36_mAd373_1 CB@36_mAd373_2 CB@36_mAd374_1 CB@36_mAd374_2 CB@36_mAd375_1 CB@36_mAd375_2 CB@36_mAd376_1 
+CB@36_mAd376_2 CB@36_mAd377_1 CB@36_mAd377_2 CB@36_mAd400_1 CB@36_mAd400_2 CB@36_mAd401_1 CB@36_mAd401_2 CB@36_mAd402_1 CB@36_mAd402_2 CB@36_mAd403_1 CB@36_mAd403_2 CB@36_mAd404_1 CB@36_mAd404_2 CB@36_mAd405_1 CB@36_mAd405_2 CB@36_mAd406_1 CB@36_mAd406_2 CB@36_mAd407_1 CB@36_mAd407_2 CB@36_mAd410_1 CB@36_mAd410_2 CB@36_mAd411_1 CB@36_mAd411_2 CB@36_mAd412_1 CB@36_mAd412_2 CB@36_mAd413_1 CB@36_mAd413_2 CB@36_mAd414_1 CB@36_mAd414_2 CB@36_mAd415_1 CB@36_mAd415_2 CB@36_mAd416_1 CB@36_mAd416_2 CB@36_mAd417_1 
+CB@36_mAd417_2 CB@36_mAd420_1 CB@36_mAd420_2 CB@36_mAd421_1 CB@36_mAd421_2 CB@36_mAd422_1 CB@36_mAd422_2 CB@36_mAd423_1 CB@36_mAd423_2 CB@36_mAd424_1 CB@36_mAd424_2 CB@36_mAd425_1 CB@36_mAd425_2 CB@36_mAd426_1 CB@36_mAd426_2 CB@36_mAd427_1 CB@36_mAd427_2 CB@36_mAd430_1 CB@36_mAd430_2 CB@36_mAd431_1 CB@36_mAd431_2 CB@36_mAd432_1 CB@36_mAd432_2 CB@36_mAd433_1 CB@36_mAd433_2 CB@36_mAd434_1 CB@36_mAd434_2 CB@36_mAd435_1 CB@36_mAd435_2 CB@36_mAd436_1 CB@36_mAd436_2 CB@36_mAd437_1 CB@36_mAd437_2 CB@36_mAd440_1 
+CB@36_mAd440_2 CB@36_mAd441_1 CB@36_mAd441_2 CB@36_mAd442_1 CB@36_mAd442_2 CB@36_mAd443_1 CB@36_mAd443_2 CB@36_mAd444_1 CB@36_mAd444_2 CB@36_mAd445_1 CB@36_mAd445_2 CB@36_mAd446_1 CB@36_mAd446_2 CB@36_mAd447_1 CB@36_mAd447_2 CB@36_mAd450_1 CB@36_mAd450_2 CB@36_mAd451_1 CB@36_mAd451_2 CB@36_mAd452_1 CB@36_mAd452_2 CB@36_mAd453_1 CB@36_mAd453_2 CB@36_mAd454_1 CB@36_mAd454_2 CB@36_mAd455_1 CB@36_mAd455_2 CB@36_mAd456_1 CB@36_mAd456_2 CB@36_mAd457_1 CB@36_mAd457_2 CB@36_mAd460_1 CB@36_mAd460_2 CB@36_mAd466_1 
+CB@36_mAd466_2 CB@36_mAd467_1 CB@36_mAd467_2 CB@36_mAd500_1 CB@36_mAd500_2 CB@36_mAd501_1 CB@36_mAd501_2 CB@36_mAd502_1 CB@36_mAd502_2 CB@36_mAd508_1 CB@36_mAd508_2 CB@36_mAd509_1 CB@36_mAd509_2 CB@36_mAd512_1 CB@36_mAd512_2 CB@36_mAd513_1 CB@36_mAd513_2 CB@36_mAd514_1 CB@36_mAd514_2 CB@36_mAd515_1 CB@36_mAd515_2 CB@36_mAd516_1 CB@36_mAd516_2 CB@36_mAd517_1 CB@36_mAd517_2 CB@36_mAd520_1 CB@36_mAd520_2 CB@36_mAd521_1 CB@36_mAd521_2 CB@36_mAd522_1 CB@36_mAd522_2 CB@36_mAd523_1 CB@36_mAd523_2 CB@36_mAd524_1 
+CB@36_mAd524_2 CB@36_mAd525_1 CB@36_mAd525_2 CB@36_mAd526_1 CB@36_mAd526_2 CB@36_mAd527_1 CB@36_mAd527_2 CB@36_mAd530_1 CB@36_mAd530_2 CB@36_mAd531_1 CB@36_mAd531_2 CB@36_mAd532_1 CB@36_mAd532_2 CB@36_mAd533_1 CB@36_mAd533_2 CB@36_mAd534_1 CB@36_mAd534_2 CB@36_mAd535_1 CB@36_mAd535_2 CB@36_mAd536_1 CB@36_mAd536_2 CB@36_mAd537_1 CB@36_mAd537_2 CB@36_mAd540_1 CB@36_mAd540_2 CB@36_mAd541_1 CB@36_mAd541_2 CB@36_mAd542_1 CB@36_mAd542_2 CB@36_mAd543_1 CB@36_mAd543_2 CB@36_mAd544_1 CB@36_mAd544_2 CB@36_mAd545_1 
+CB@36_mAd545_2 CB@36_mAd546_1 CB@36_mAd546_2 CB@36_mAd547_1 CB@36_mAd547_2 CB@36_mAd550_1 CB@36_mAd550_2 CB@36_mAd551_1 CB@36_mAd551_2 CB@36_mAd552_1 CB@36_mAd552_2 CB@36_mAd553_1 CB@36_mAd553_2 CB@36_mAd554_1 CB@36_mAd554_2 CB@36_mAd555_1 CB@36_mAd555_2 CB@36_mAd556_1 CB@36_mAd556_2 CB@36_mAd557_1 CB@36_mAd557_2 CB@36_mAd560_1 CB@36_mAd560_2 CB@36_mAd561_1 CB@36_mAd561_2 CB@36_mAd562_1 CB@36_mAd562_2 CB@36_mAd563_1 CB@36_mAd563_2 CB@36_mAd564_1 CB@36_mAd564_2 CB@36_mAd565_1 CB@36_mAd565_2 CB@36_mAd566_1 
+CB@36_mAd566_2 CB@36_mAd567_1 CB@36_mAd567_2 CB@36_mAd570_1 CB@36_mAd570_2 CB@36_mAd571_1 CB@36_mAd571_2 CB@36_mAd572_1 CB@36_mAd572_2 CB@36_mAd573_1 CB@36_mAd573_2 CB@36_mAd575_1 CB@36_mAd575_2 CB@36_mAd576_1 CB@36_mAd576_2 CB@36_mAd577_1 CB@36_mAd577_2 CB@36_mAd600_1 CB@36_mAd600_2 CB@36_mAd601_1 CB@36_mAd601_2 CB@36_mAd602_1 CB@36_mAd602_2 CB@36_mAd604_1 CB@36_mAd604_2 CB@36_mAd605_1 CB@36_mAd605_2 CB@36_mAd606_1 CB@36_mAd606_2 CB@36_mAd607_1 CB@36_mAd607_2 CB@36_mAd610_1 CB@36_mAd610_2 CB@36_mAd611_1 
+CB@36_mAd611_2 CB@36_mAd612_1 CB@36_mAd612_2 CB@36_mAd613_1 CB@36_mAd613_2 CB@36_mAd614_1 CB@36_mAd614_2 CB@36_mAd615_1 CB@36_mAd615_2 CB@36_mAd616_1 CB@36_mAd616_2 CB@36_mAd617_1 CB@36_mAd617_2 CB@36_mAd620_1 CB@36_mAd620_2 CB@36_mAd621_1 CB@36_mAd621_2 CB@36_mAd622_1 CB@36_mAd622_2 CB@36_mAd623_1 CB@36_mAd623_2 CB@36_mAd624_1 CB@36_mAd624_2 CB@36_mAd625_1 CB@36_mAd625_2 CB@36_mAd626_1 CB@36_mAd626_2 CB@36_mAd627_1 CB@36_mAd627_2 CB@36_mAd630_1 CB@36_mAd630_2 CB@36_mAd631_1 CB@36_mAd631_2 CB@36_mAd632_1 
+CB@36_mAd632_2 CB@36_mAd633_1 CB@36_mAd633_2 CB@36_mAd634_1 CB@36_mAd634_2 CB@36_mAd635_1 CB@36_mAd635_2 CB@36_mAd636_1 CB@36_mAd636_2 CB@36_mAd637_1 CB@36_mAd637_2 CB@36_mAd640_1 CB@36_mAd640_2 CB@36_mAd641_1 CB@36_mAd641_2 CB@36_mAd642_1 CB@36_mAd642_2 CB@36_mAd643_1 CB@36_mAd643_2 CB@36_mAd644_1 CB@36_mAd644_2 CB@36_mAd645_1 CB@36_mAd645_2 CB@36_mAd646_1 CB@36_mAd646_2 CB@36_mAd647_1 CB@36_mAd647_2 CB@36_mAd650_1 CB@36_mAd650_2 CB@36_mAd651_1 CB@36_mAd651_2 CB@36_mAd652_1 CB@36_mAd652_2 CB@36_mAd653_1 
+CB@36_mAd653_2 CB@36_mAd654_1 CB@36_mAd654_2 CB@36_mAd655_1 CB@36_mAd655_2 CB@36_mAd656_1 CB@36_mAd656_2 CB@36_mAd657_1 CB@36_mAd657_2 CB@36_mAd660_1 CB@36_mAd660_2 CB@36_mAd661_1 CB@36_mAd661_2 CB@36_mAd662_1 CB@36_mAd662_2 CB@36_mAd663_1 CB@36_mAd663_2 CB@36_mAd664_1 CB@36_mAd664_2 CB@36_mAd665_1 CB@36_mAd665_2 CB@36_mAd666_1 CB@36_mAd666_2 CB@36_mAd667_1 CB@36_mAd667_2 CB@36_mAd675_1 CB@36_mAd675_2 CB@36_mAd676_1 CB@36_mAd676_2 CB@36_mAd677_1 CB@36_mAd677_2 CB@36_mAd700_1 CB@36_mAd700_2 CB@36_mAd710_1 
+CB@36_mAd710_2 CB@36_mAd711_1 CB@36_mAd711_2 CB@36_mAd717_1 CB@36_mAd717_2 CB@36_mAd720_1 CB@36_mAd720_2 CB@36_mAd721_1 CB@36_mAd721_2 CB@36_mAd722_1 CB@36_mAd722_2 CB@36_mAd723_1 CB@36_mAd723_2 CB@36_mAd724_1 CB@36_mAd724_2 CB@36_mAd725_1 CB@36_mAd725_2 CB@36_mAd726_1 CB@36_mAd726_2 CB@36_mAd727_1 CB@36_mAd727_2 CB@36_mAd730_1 CB@36_mAd730_2 CB@36_mAd731_1 CB@36_mAd731_2 CB@36_mAd732_1 CB@36_mAd732_2 CB@36_mAd733_1 CB@36_mAd733_2 CB@36_mAd734_1 CB@36_mAd734_2 CB@36_mAd735_1 CB@36_mAd735_2 CB@36_mAd736_1 
+CB@36_mAd736_2 CB@36_mAd737_1 CB@36_mAd737_2 CB@36_mAd740_1 CB@36_mAd740_2 CB@36_mAd741_1 CB@36_mAd741_2 CB@36_mAd742_1 CB@36_mAd742_2 CB@36_mAd743_1 CB@36_mAd743_2 CB@36_mAd744_1 CB@36_mAd744_2 CB@36_mAd745_1 CB@36_mAd745_2 CB@36_mAd746_1 CB@36_mAd746_2 CB@36_mAd747_1 CB@36_mAd747_2 CB@36_mAd750_1 CB@36_mAd750_2 CB@36_mAd751_1 CB@36_mAd751_2 CB@36_mAd752_1 CB@36_mAd752_2 CB@36_mAd753_1 CB@36_mAd753_2 CB@36_mAd754_1 CB@36_mAd754_2 CB@36_mAd755_1 CB@36_mAd755_2 CB@36_mAd756_1 CB@36_mAd756_2 CB@36_mAd757_1 
+CB@36_mAd757_2 CB@36_mAd760_1 CB@36_mAd760_2 CB@36_mAd761_1 CB@36_mAd761_2 CB@36_mAd762_1 CB@36_mAd762_2 CB@36_mAd763_1 CB@36_mAd763_2 CB@36_mAd764_1 CB@36_mAd764_2 CB@36_mAd765_1 CB@36_mAd765_2 CB@36_mAd766_1 CB@36_mAd766_2 CB@36_mAd767_1 CB@36_mAd767_2 CB@36_mAd771_1 CB@36_mAd771_2 CB@36_mAd772_1 CB@36_mAd772_2 CB@36_mAd773_1 CB@36_mAd773_2 CB@36_mAd774_1 CB@36_mAd774_2 CB@36_mAd775_1 CB@36_mAd775_2 CB@36_mAd776_1 CB@36_mAd776_2 CB@36_mAd777_1 CB@36_mAd777_2 CB@36_X0 CB@36_X1 CB@36_X10 CB@36_X11 
+CB@36_X12 CB@36_X13 CB@36_X2 CB@36_X3 CB@36_X4 CB@36_X5 CB@36_X6 CB@36_X7 CB@36_X8 CB@36_X9 CB@36_Y1 CB@36_Y10 CB@36_Y11 CB@36_Y12 CB@36_Y2 CB@36_Y3 CB@36_Y4 CB@36_Y5 CB@36_Y6 CB@36_Y7 CB@36_Y8 CB@36_Y9 CB@36_Z1 CB@36_Z10 CB@36_Z11 CB@36_Z12 CB@36_Z2 CB@36_Z3 CB@36_Z4 CB@36_Z5 CB@36_Z6 CB@36_Z7 CB@36_Z8 CB@36_Z9 _5400TP094__CB
XCB@37 CB@37_K0 CB@37_K1 CB@37_K10 CB@37_K11 CB@37_K12 CB@37_K13 CB@37_K2 CB@37_K3 CB@37_K4 CB@37_K5 CB@37_K6 CB@37_K7 CB@37_K8 CB@37_K9 CB@37_mAd000_1 CB@37_mAd000_2 CB@37_mAd001_1 CB@37_mAd001_2 CB@37_mAd002_1 CB@37_mAd002_2 CB@37_mAd003_1 CB@37_mAd003_2 CB@37_mAd004_1 CB@37_mAd004_2 CB@37_mAd005_1 CB@37_mAd005_2 CB@37_mAd006_1 CB@37_mAd006_2 CB@37_mAd007_1 CB@37_mAd007_2 CB@37_mAd010_1 CB@37_mAd010_2 CB@37_mAd011_1 CB@37_mAd011_2 CB@37_mAd012_1 CB@37_mAd012_2 CB@37_mAd013_1 CB@37_mAd013_2 CB@37_mAd014_1 
+CB@37_mAd014_2 CB@37_mAd015_1 CB@37_mAd015_2 CB@37_mAd016_1 CB@37_mAd016_2 CB@37_mAd017_1 CB@37_mAd017_2 CB@37_mAd020_1 CB@37_mAd020_2 CB@37_mAd021_1 CB@37_mAd021_2 CB@37_mAd022_1 CB@37_mAd022_2 CB@37_mAd023_1 CB@37_mAd023_2 CB@37_mAd024_1 CB@37_mAd024_2 CB@37_mAd025_1 CB@37_mAd025_2 CB@37_mAd026_1 CB@37_mAd026_2 CB@37_mAd027_1 CB@37_mAd027_2 CB@37_mAd030_1 CB@37_mAd030_2 CB@37_mAd031_1 CB@37_mAd031_2 CB@37_mAd032_1 CB@37_mAd032_2 CB@37_mAd033_1 CB@37_mAd033_2 CB@37_mAd034_1 CB@37_mAd034_2 CB@37_mAd035_1 
+CB@37_mAd035_2 CB@37_mAd036_1 CB@37_mAd036_2 CB@37_mAd037_1 CB@37_mAd037_2 CB@37_mAd040_1 CB@37_mAd040_2 CB@37_mAd041_1 CB@37_mAd041_2 CB@37_mAd042_1 CB@37_mAd042_2 CB@37_mAd043_1 CB@37_mAd043_2 CB@37_mAd044_1 CB@37_mAd044_2 CB@37_mAd045_1 CB@37_mAd045_2 CB@37_mAd046_1 CB@37_mAd046_2 CB@37_mAd047_1 CB@37_mAd047_2 CB@37_mAd050_1 CB@37_mAd050_2 CB@37_mAd051_1 CB@37_mAd051_2 CB@37_mAd052_1 CB@37_mAd052_2 CB@37_mAd053_1 CB@37_mAd053_2 CB@37_mAd054_1 CB@37_mAd054_2 CB@37_mAd055_1 CB@37_mAd055_2 CB@37_mAd056_1 
+CB@37_mAd056_2 CB@37_mAd057_1 CB@37_mAd057_2 CB@37_mAd060_1 CB@37_mAd060_2 CB@37_mAd066_1 CB@37_mAd066_2 CB@37_mAd067_1 CB@37_mAd067_2 CB@37_mAd100_1 CB@37_mAd100_2 CB@37_mAd101_1 CB@37_mAd101_2 CB@37_mAd102_1 CB@37_mAd102_2 CB@37_mAd110_1 CB@37_mAd110_2 CB@37_mAd111_1 CB@37_mAd111_2 CB@37_mAd112_1 CB@37_mAd112_2 CB@37_mAd113_1 CB@37_mAd113_2 CB@37_mAd114_1 CB@37_mAd114_2 CB@37_mAd115_1 CB@37_mAd115_2 CB@37_mAd116_1 CB@37_mAd116_2 CB@37_mAd117_1 CB@37_mAd117_2 CB@37_mAd120_1 CB@37_mAd120_2 CB@37_mAd121_1 
+CB@37_mAd121_2 CB@37_mAd122_1 CB@37_mAd122_2 CB@37_mAd123_1 CB@37_mAd123_2 CB@37_mAd124_1 CB@37_mAd124_2 CB@37_mAd125_1 CB@37_mAd125_2 CB@37_mAd126_1 CB@37_mAd126_2 CB@37_mAd127_1 CB@37_mAd127_2 CB@37_mAd130_1 CB@37_mAd130_2 CB@37_mAd131_1 CB@37_mAd131_2 CB@37_mAd132_1 CB@37_mAd132_2 CB@37_mAd133_1 CB@37_mAd133_2 CB@37_mAd134_1 CB@37_mAd134_2 CB@37_mAd135_1 CB@37_mAd135_2 CB@37_mAd136_1 CB@37_mAd136_2 CB@37_mAd137_1 CB@37_mAd137_2 CB@37_mAd140_1 CB@37_mAd140_2 CB@37_mAd141_1 CB@37_mAd141_2 CB@37_mAd142_1 
+CB@37_mAd142_2 CB@37_mAd143_1 CB@37_mAd143_2 CB@37_mAd144_1 CB@37_mAd144_2 CB@37_mAd145_1 CB@37_mAd145_2 CB@37_mAd146_1 CB@37_mAd146_2 CB@37_mAd147_1 CB@37_mAd147_2 CB@37_mAd150_1 CB@37_mAd150_2 CB@37_mAd151_1 CB@37_mAd151_2 CB@37_mAd152_1 CB@37_mAd152_2 CB@37_mAd153_1 CB@37_mAd153_2 CB@37_mAd154_1 CB@37_mAd154_2 CB@37_mAd155_1 CB@37_mAd155_2 CB@37_mAd156_1 CB@37_mAd156_2 CB@37_mAd157_1 CB@37_mAd157_2 CB@37_mAd160_1 CB@37_mAd160_2 CB@37_mAd161_1 CB@37_mAd161_2 CB@37_mAd162_1 CB@37_mAd162_2 CB@37_mAd163_1 
+CB@37_mAd163_2 CB@37_mAd164_1 CB@37_mAd164_2 CB@37_mAd165_1 CB@37_mAd165_2 CB@37_mAd166_1 CB@37_mAd166_2 CB@37_mAd167_1 CB@37_mAd167_2 CB@37_mAd170_1 CB@37_mAd170_2 CB@37_mAd171_1 CB@37_mAd171_2 CB@37_mAd172_1 CB@37_mAd172_2 CB@37_mAd173_1 CB@37_mAd173_2 CB@37_mAd175_1 CB@37_mAd175_2 CB@37_mAd176_1 CB@37_mAd176_2 CB@37_mAd177_1 CB@37_mAd177_2 CB@37_mAd200_1 CB@37_mAd200_2 CB@37_mAd201_1 CB@37_mAd201_2 CB@37_mAd202_1 CB@37_mAd202_2 CB@37_mAd204_1 CB@37_mAd204_2 CB@37_mAd205_1 CB@37_mAd205_2 CB@37_mAd206_1 
+CB@37_mAd206_2 CB@37_mAd207_1 CB@37_mAd207_2 CB@37_mAd210_1 CB@37_mAd210_2 CB@37_mAd211_1 CB@37_mAd211_2 CB@37_mAd212_1 CB@37_mAd212_2 CB@37_mAd213_1 CB@37_mAd213_2 CB@37_mAd214_1 CB@37_mAd214_2 CB@37_mAd215_1 CB@37_mAd215_2 CB@37_mAd216_1 CB@37_mAd216_2 CB@37_mAd217_1 CB@37_mAd217_2 CB@37_mAd220_1 CB@37_mAd220_2 CB@37_mAd221_1 CB@37_mAd221_2 CB@37_mAd222_1 CB@37_mAd222_2 CB@37_mAd223_1 CB@37_mAd223_2 CB@37_mAd224_1 CB@37_mAd224_2 CB@37_mAd225_1 CB@37_mAd225_2 CB@37_mAd226_1 CB@37_mAd226_2 CB@37_mAd227_1 
+CB@37_mAd227_2 CB@37_mAd230_1 CB@37_mAd230_2 CB@37_mAd231_1 CB@37_mAd231_2 CB@37_mAd232_1 CB@37_mAd232_2 CB@37_mAd233_1 CB@37_mAd233_2 CB@37_mAd234_1 CB@37_mAd234_2 CB@37_mAd235_1 CB@37_mAd235_2 CB@37_mAd236_1 CB@37_mAd236_2 CB@37_mAd237_1 CB@37_mAd237_2 CB@37_mAd240_1 CB@37_mAd240_2 CB@37_mAd241_1 CB@37_mAd241_2 CB@37_mAd242_1 CB@37_mAd242_2 CB@37_mAd243_1 CB@37_mAd243_2 CB@37_mAd244_1 CB@37_mAd244_2 CB@37_mAd245_1 CB@37_mAd245_2 CB@37_mAd246_1 CB@37_mAd246_2 CB@37_mAd247_1 CB@37_mAd247_2 CB@37_mAd250_1 
+CB@37_mAd250_2 CB@37_mAd251_1 CB@37_mAd251_2 CB@37_mAd252_1 CB@37_mAd252_2 CB@37_mAd253_1 CB@37_mAd253_2 CB@37_mAd254_1 CB@37_mAd254_2 CB@37_mAd255_1 CB@37_mAd255_2 CB@37_mAd256_1 CB@37_mAd256_2 CB@37_mAd257_1 CB@37_mAd257_2 CB@37_mAd260_1 CB@37_mAd260_2 CB@37_mAd261_1 CB@37_mAd261_2 CB@37_mAd262_1 CB@37_mAd262_2 CB@37_mAd263_1 CB@37_mAd263_2 CB@37_mAd264_1 CB@37_mAd264_2 CB@37_mAd265_1 CB@37_mAd265_2 CB@37_mAd266_1 CB@37_mAd266_2 CB@37_mAd267_1 CB@37_mAd267_2 CB@37_mAd275_1 CB@37_mAd275_2 CB@37_mAd276_1 
+CB@37_mAd276_2 CB@37_mAd277_1 CB@37_mAd277_2 CB@37_mAd300_1 CB@37_mAd300_2 CB@37_mAd310_1 CB@37_mAd310_2 CB@37_mAd311_1 CB@37_mAd311_2 CB@37_mAd317_1 CB@37_mAd317_2 CB@37_mAd320_1 CB@37_mAd320_2 CB@37_mAd321_1 CB@37_mAd321_2 CB@37_mAd322_1 CB@37_mAd322_2 CB@37_mAd323_1 CB@37_mAd323_2 CB@37_mAd324_1 CB@37_mAd324_2 CB@37_mAd325_1 CB@37_mAd325_2 CB@37_mAd326_1 CB@37_mAd326_2 CB@37_mAd327_1 CB@37_mAd327_2 CB@37_mAd330_1 CB@37_mAd330_2 CB@37_mAd331_1 CB@37_mAd331_2 CB@37_mAd332_1 CB@37_mAd332_2 CB@37_mAd333_1 
+CB@37_mAd333_2 CB@37_mAd334_1 CB@37_mAd334_2 CB@37_mAd335_1 CB@37_mAd335_2 CB@37_mAd336_1 CB@37_mAd336_2 CB@37_mAd337_1 CB@37_mAd337_2 CB@37_mAd340_1 CB@37_mAd340_2 CB@37_mAd341_1 CB@37_mAd341_2 CB@37_mAd342_1 CB@37_mAd342_2 CB@37_mAd343_1 CB@37_mAd343_2 CB@37_mAd344_1 CB@37_mAd344_2 CB@37_mAd345_1 CB@37_mAd345_2 CB@37_mAd346_1 CB@37_mAd346_2 CB@37_mAd347_1 CB@37_mAd347_2 CB@37_mAd350_1 CB@37_mAd350_2 CB@37_mAd351_1 CB@37_mAd351_2 CB@37_mAd352_1 CB@37_mAd352_2 CB@37_mAd353_1 CB@37_mAd353_2 CB@37_mAd354_1 
+CB@37_mAd354_2 CB@37_mAd355_1 CB@37_mAd355_2 CB@37_mAd356_1 CB@37_mAd356_2 CB@37_mAd357_1 CB@37_mAd357_2 CB@37_mAd360_1 CB@37_mAd360_2 CB@37_mAd361_1 CB@37_mAd361_2 CB@37_mAd362_1 CB@37_mAd362_2 CB@37_mAd363_1 CB@37_mAd363_2 CB@37_mAd364_1 CB@37_mAd364_2 CB@37_mAd365_1 CB@37_mAd365_2 CB@37_mAd366_1 CB@37_mAd366_2 CB@37_mAd367_1 CB@37_mAd367_2 CB@37_mAd371_1 CB@37_mAd371_2 CB@37_mAd372_1 CB@37_mAd372_2 CB@37_mAd373_1 CB@37_mAd373_2 CB@37_mAd374_1 CB@37_mAd374_2 CB@37_mAd375_1 CB@37_mAd375_2 CB@37_mAd376_1 
+CB@37_mAd376_2 CB@37_mAd377_1 CB@37_mAd377_2 CB@37_mAd400_1 CB@37_mAd400_2 CB@37_mAd401_1 CB@37_mAd401_2 CB@37_mAd402_1 CB@37_mAd402_2 CB@37_mAd403_1 CB@37_mAd403_2 CB@37_mAd404_1 CB@37_mAd404_2 CB@37_mAd405_1 CB@37_mAd405_2 CB@37_mAd406_1 CB@37_mAd406_2 CB@37_mAd407_1 CB@37_mAd407_2 CB@37_mAd410_1 CB@37_mAd410_2 CB@37_mAd411_1 CB@37_mAd411_2 CB@37_mAd412_1 CB@37_mAd412_2 CB@37_mAd413_1 CB@37_mAd413_2 CB@37_mAd414_1 CB@37_mAd414_2 CB@37_mAd415_1 CB@37_mAd415_2 CB@37_mAd416_1 CB@37_mAd416_2 CB@37_mAd417_1 
+CB@37_mAd417_2 CB@37_mAd420_1 CB@37_mAd420_2 CB@37_mAd421_1 CB@37_mAd421_2 CB@37_mAd422_1 CB@37_mAd422_2 CB@37_mAd423_1 CB@37_mAd423_2 CB@37_mAd424_1 CB@37_mAd424_2 CB@37_mAd425_1 CB@37_mAd425_2 CB@37_mAd426_1 CB@37_mAd426_2 CB@37_mAd427_1 CB@37_mAd427_2 CB@37_mAd430_1 CB@37_mAd430_2 CB@37_mAd431_1 CB@37_mAd431_2 CB@37_mAd432_1 CB@37_mAd432_2 CB@37_mAd433_1 CB@37_mAd433_2 CB@37_mAd434_1 CB@37_mAd434_2 CB@37_mAd435_1 CB@37_mAd435_2 CB@37_mAd436_1 CB@37_mAd436_2 CB@37_mAd437_1 CB@37_mAd437_2 CB@37_mAd440_1 
+CB@37_mAd440_2 CB@37_mAd441_1 CB@37_mAd441_2 CB@37_mAd442_1 CB@37_mAd442_2 CB@37_mAd443_1 CB@37_mAd443_2 CB@37_mAd444_1 CB@37_mAd444_2 CB@37_mAd445_1 CB@37_mAd445_2 CB@37_mAd446_1 CB@37_mAd446_2 CB@37_mAd447_1 CB@37_mAd447_2 CB@37_mAd450_1 CB@37_mAd450_2 CB@37_mAd451_1 CB@37_mAd451_2 CB@37_mAd452_1 CB@37_mAd452_2 CB@37_mAd453_1 CB@37_mAd453_2 CB@37_mAd454_1 CB@37_mAd454_2 CB@37_mAd455_1 CB@37_mAd455_2 CB@37_mAd456_1 CB@37_mAd456_2 CB@37_mAd457_1 CB@37_mAd457_2 CB@37_mAd460_1 CB@37_mAd460_2 CB@37_mAd466_1 
+CB@37_mAd466_2 CB@37_mAd467_1 CB@37_mAd467_2 CB@37_mAd500_1 CB@37_mAd500_2 CB@37_mAd501_1 CB@37_mAd501_2 CB@37_mAd502_1 CB@37_mAd502_2 CB@37_mAd508_1 CB@37_mAd508_2 CB@37_mAd509_1 CB@37_mAd509_2 CB@37_mAd512_1 CB@37_mAd512_2 CB@37_mAd513_1 CB@37_mAd513_2 CB@37_mAd514_1 CB@37_mAd514_2 CB@37_mAd515_1 CB@37_mAd515_2 CB@37_mAd516_1 CB@37_mAd516_2 CB@37_mAd517_1 CB@37_mAd517_2 CB@37_mAd520_1 CB@37_mAd520_2 CB@37_mAd521_1 CB@37_mAd521_2 CB@37_mAd522_1 CB@37_mAd522_2 CB@37_mAd523_1 CB@37_mAd523_2 CB@37_mAd524_1 
+CB@37_mAd524_2 CB@37_mAd525_1 CB@37_mAd525_2 CB@37_mAd526_1 CB@37_mAd526_2 CB@37_mAd527_1 CB@37_mAd527_2 CB@37_mAd530_1 CB@37_mAd530_2 CB@37_mAd531_1 CB@37_mAd531_2 CB@37_mAd532_1 CB@37_mAd532_2 CB@37_mAd533_1 CB@37_mAd533_2 CB@37_mAd534_1 CB@37_mAd534_2 CB@37_mAd535_1 CB@37_mAd535_2 CB@37_mAd536_1 CB@37_mAd536_2 CB@37_mAd537_1 CB@37_mAd537_2 CB@37_mAd540_1 CB@37_mAd540_2 CB@37_mAd541_1 CB@37_mAd541_2 CB@37_mAd542_1 CB@37_mAd542_2 CB@37_mAd543_1 CB@37_mAd543_2 CB@37_mAd544_1 CB@37_mAd544_2 CB@37_mAd545_1 
+CB@37_mAd545_2 CB@37_mAd546_1 CB@37_mAd546_2 CB@37_mAd547_1 CB@37_mAd547_2 CB@37_mAd550_1 CB@37_mAd550_2 CB@37_mAd551_1 CB@37_mAd551_2 CB@37_mAd552_1 CB@37_mAd552_2 CB@37_mAd553_1 CB@37_mAd553_2 CB@37_mAd554_1 CB@37_mAd554_2 CB@37_mAd555_1 CB@37_mAd555_2 CB@37_mAd556_1 CB@37_mAd556_2 CB@37_mAd557_1 CB@37_mAd557_2 CB@37_mAd560_1 CB@37_mAd560_2 CB@37_mAd561_1 CB@37_mAd561_2 CB@37_mAd562_1 CB@37_mAd562_2 CB@37_mAd563_1 CB@37_mAd563_2 CB@37_mAd564_1 CB@37_mAd564_2 CB@37_mAd565_1 CB@37_mAd565_2 CB@37_mAd566_1 
+CB@37_mAd566_2 CB@37_mAd567_1 CB@37_mAd567_2 CB@37_mAd570_1 CB@37_mAd570_2 CB@37_mAd571_1 CB@37_mAd571_2 CB@37_mAd572_1 CB@37_mAd572_2 CB@37_mAd573_1 CB@37_mAd573_2 CB@37_mAd575_1 CB@37_mAd575_2 CB@37_mAd576_1 CB@37_mAd576_2 CB@37_mAd577_1 CB@37_mAd577_2 CB@37_mAd600_1 CB@37_mAd600_2 CB@37_mAd601_1 CB@37_mAd601_2 CB@37_mAd602_1 CB@37_mAd602_2 CB@37_mAd604_1 CB@37_mAd604_2 CB@37_mAd605_1 CB@37_mAd605_2 CB@37_mAd606_1 CB@37_mAd606_2 CB@37_mAd607_1 CB@37_mAd607_2 CB@37_mAd610_1 CB@37_mAd610_2 CB@37_mAd611_1 
+CB@37_mAd611_2 CB@37_mAd612_1 CB@37_mAd612_2 CB@37_mAd613_1 CB@37_mAd613_2 CB@37_mAd614_1 CB@37_mAd614_2 CB@37_mAd615_1 CB@37_mAd615_2 CB@37_mAd616_1 CB@37_mAd616_2 CB@37_mAd617_1 CB@37_mAd617_2 CB@37_mAd620_1 CB@37_mAd620_2 CB@37_mAd621_1 CB@37_mAd621_2 CB@37_mAd622_1 CB@37_mAd622_2 CB@37_mAd623_1 CB@37_mAd623_2 CB@37_mAd624_1 CB@37_mAd624_2 CB@37_mAd625_1 CB@37_mAd625_2 CB@37_mAd626_1 CB@37_mAd626_2 CB@37_mAd627_1 CB@37_mAd627_2 CB@37_mAd630_1 CB@37_mAd630_2 CB@37_mAd631_1 CB@37_mAd631_2 CB@37_mAd632_1 
+CB@37_mAd632_2 CB@37_mAd633_1 CB@37_mAd633_2 CB@37_mAd634_1 CB@37_mAd634_2 CB@37_mAd635_1 CB@37_mAd635_2 CB@37_mAd636_1 CB@37_mAd636_2 CB@37_mAd637_1 CB@37_mAd637_2 CB@37_mAd640_1 CB@37_mAd640_2 CB@37_mAd641_1 CB@37_mAd641_2 CB@37_mAd642_1 CB@37_mAd642_2 CB@37_mAd643_1 CB@37_mAd643_2 CB@37_mAd644_1 CB@37_mAd644_2 CB@37_mAd645_1 CB@37_mAd645_2 CB@37_mAd646_1 CB@37_mAd646_2 CB@37_mAd647_1 CB@37_mAd647_2 CB@37_mAd650_1 CB@37_mAd650_2 CB@37_mAd651_1 CB@37_mAd651_2 CB@37_mAd652_1 CB@37_mAd652_2 CB@37_mAd653_1 
+CB@37_mAd653_2 CB@37_mAd654_1 CB@37_mAd654_2 CB@37_mAd655_1 CB@37_mAd655_2 CB@37_mAd656_1 CB@37_mAd656_2 CB@37_mAd657_1 CB@37_mAd657_2 CB@37_mAd660_1 CB@37_mAd660_2 CB@37_mAd661_1 CB@37_mAd661_2 CB@37_mAd662_1 CB@37_mAd662_2 CB@37_mAd663_1 CB@37_mAd663_2 CB@37_mAd664_1 CB@37_mAd664_2 CB@37_mAd665_1 CB@37_mAd665_2 CB@37_mAd666_1 CB@37_mAd666_2 CB@37_mAd667_1 CB@37_mAd667_2 CB@37_mAd675_1 CB@37_mAd675_2 CB@37_mAd676_1 CB@37_mAd676_2 CB@37_mAd677_1 CB@37_mAd677_2 CB@37_mAd700_1 CB@37_mAd700_2 CB@37_mAd710_1 
+CB@37_mAd710_2 CB@37_mAd711_1 CB@37_mAd711_2 CB@37_mAd717_1 CB@37_mAd717_2 CB@37_mAd720_1 CB@37_mAd720_2 CB@37_mAd721_1 CB@37_mAd721_2 CB@37_mAd722_1 CB@37_mAd722_2 CB@37_mAd723_1 CB@37_mAd723_2 CB@37_mAd724_1 CB@37_mAd724_2 CB@37_mAd725_1 CB@37_mAd725_2 CB@37_mAd726_1 CB@37_mAd726_2 CB@37_mAd727_1 CB@37_mAd727_2 CB@37_mAd730_1 CB@37_mAd730_2 CB@37_mAd731_1 CB@37_mAd731_2 CB@37_mAd732_1 CB@37_mAd732_2 CB@37_mAd733_1 CB@37_mAd733_2 CB@37_mAd734_1 CB@37_mAd734_2 CB@37_mAd735_1 CB@37_mAd735_2 CB@37_mAd736_1 
+CB@37_mAd736_2 CB@37_mAd737_1 CB@37_mAd737_2 CB@37_mAd740_1 CB@37_mAd740_2 CB@37_mAd741_1 CB@37_mAd741_2 CB@37_mAd742_1 CB@37_mAd742_2 CB@37_mAd743_1 CB@37_mAd743_2 CB@37_mAd744_1 CB@37_mAd744_2 CB@37_mAd745_1 CB@37_mAd745_2 CB@37_mAd746_1 CB@37_mAd746_2 CB@37_mAd747_1 CB@37_mAd747_2 CB@37_mAd750_1 CB@37_mAd750_2 CB@37_mAd751_1 CB@37_mAd751_2 CB@37_mAd752_1 CB@37_mAd752_2 CB@37_mAd753_1 CB@37_mAd753_2 CB@37_mAd754_1 CB@37_mAd754_2 CB@37_mAd755_1 CB@37_mAd755_2 CB@37_mAd756_1 CB@37_mAd756_2 CB@37_mAd757_1 
+CB@37_mAd757_2 CB@37_mAd760_1 CB@37_mAd760_2 CB@37_mAd761_1 CB@37_mAd761_2 CB@37_mAd762_1 CB@37_mAd762_2 CB@37_mAd763_1 CB@37_mAd763_2 CB@37_mAd764_1 CB@37_mAd764_2 CB@37_mAd765_1 CB@37_mAd765_2 CB@37_mAd766_1 CB@37_mAd766_2 CB@37_mAd767_1 CB@37_mAd767_2 CB@37_mAd771_1 CB@37_mAd771_2 CB@37_mAd772_1 CB@37_mAd772_2 CB@37_mAd773_1 CB@37_mAd773_2 CB@37_mAd774_1 CB@37_mAd774_2 CB@37_mAd775_1 CB@37_mAd775_2 CB@37_mAd776_1 CB@37_mAd776_2 CB@37_mAd777_1 CB@37_mAd777_2 CB@37_X0 CB@37_X1 CB@37_X10 CB@37_X11 
+CB@37_X12 CB@37_X13 CB@37_X2 CB@37_X3 CB@37_X4 CB@37_X5 CB@37_X6 CB@37_X7 CB@37_X8 CB@37_X9 CB@37_Y1 CB@37_Y10 CB@37_Y11 CB@37_Y12 CB@37_Y2 CB@37_Y3 CB@37_Y4 CB@37_Y5 CB@37_Y6 CB@37_Y7 CB@37_Y8 CB@37_Y9 CB@37_Z1 CB@37_Z10 CB@37_Z11 CB@37_Z12 CB@37_Z2 CB@37_Z3 CB@37_Z4 CB@37_Z5 CB@37_Z6 CB@37_Z7 CB@37_Z8 CB@37_Z9 _5400TP094__CB
XCB@38 CB@38_K0 CB@38_K1 CB@38_K10 CB@38_K11 CB@38_K12 CB@38_K13 CB@38_K2 CB@38_K3 CB@38_K4 CB@38_K5 CB@38_K6 CB@38_K7 CB@38_K8 CB@38_K9 CB@38_mAd000_1 CB@38_mAd000_2 CB@38_mAd001_1 CB@38_mAd001_2 CB@38_mAd002_1 CB@38_mAd002_2 CB@38_mAd003_1 CB@38_mAd003_2 CB@38_mAd004_1 CB@38_mAd004_2 CB@38_mAd005_1 CB@38_mAd005_2 CB@38_mAd006_1 CB@38_mAd006_2 CB@38_mAd007_1 CB@38_mAd007_2 CB@38_mAd010_1 CB@38_mAd010_2 CB@38_mAd011_1 CB@38_mAd011_2 CB@38_mAd012_1 CB@38_mAd012_2 CB@38_mAd013_1 CB@38_mAd013_2 CB@38_mAd014_1 
+CB@38_mAd014_2 CB@38_mAd015_1 CB@38_mAd015_2 CB@38_mAd016_1 CB@38_mAd016_2 CB@38_mAd017_1 CB@38_mAd017_2 CB@38_mAd020_1 CB@38_mAd020_2 CB@38_mAd021_1 CB@38_mAd021_2 CB@38_mAd022_1 CB@38_mAd022_2 CB@38_mAd023_1 CB@38_mAd023_2 CB@38_mAd024_1 CB@38_mAd024_2 CB@38_mAd025_1 CB@38_mAd025_2 CB@38_mAd026_1 CB@38_mAd026_2 CB@38_mAd027_1 CB@38_mAd027_2 CB@38_mAd030_1 CB@38_mAd030_2 CB@38_mAd031_1 CB@38_mAd031_2 CB@38_mAd032_1 CB@38_mAd032_2 CB@38_mAd033_1 CB@38_mAd033_2 CB@38_mAd034_1 CB@38_mAd034_2 CB@38_mAd035_1 
+CB@38_mAd035_2 CB@38_mAd036_1 CB@38_mAd036_2 CB@38_mAd037_1 CB@38_mAd037_2 CB@38_mAd040_1 CB@38_mAd040_2 CB@38_mAd041_1 CB@38_mAd041_2 CB@38_mAd042_1 CB@38_mAd042_2 CB@38_mAd043_1 CB@38_mAd043_2 CB@38_mAd044_1 CB@38_mAd044_2 CB@38_mAd045_1 CB@38_mAd045_2 CB@38_mAd046_1 CB@38_mAd046_2 CB@38_mAd047_1 CB@38_mAd047_2 CB@38_mAd050_1 CB@38_mAd050_2 CB@38_mAd051_1 CB@38_mAd051_2 CB@38_mAd052_1 CB@38_mAd052_2 CB@38_mAd053_1 CB@38_mAd053_2 CB@38_mAd054_1 CB@38_mAd054_2 CB@38_mAd055_1 CB@38_mAd055_2 CB@38_mAd056_1 
+CB@38_mAd056_2 CB@38_mAd057_1 CB@38_mAd057_2 CB@38_mAd060_1 CB@38_mAd060_2 CB@38_mAd066_1 CB@38_mAd066_2 CB@38_mAd067_1 CB@38_mAd067_2 CB@38_mAd100_1 CB@38_mAd100_2 CB@38_mAd101_1 CB@38_mAd101_2 CB@38_mAd102_1 CB@38_mAd102_2 CB@38_mAd110_1 CB@38_mAd110_2 CB@38_mAd111_1 CB@38_mAd111_2 CB@38_mAd112_1 CB@38_mAd112_2 CB@38_mAd113_1 CB@38_mAd113_2 CB@38_mAd114_1 CB@38_mAd114_2 CB@38_mAd115_1 CB@38_mAd115_2 CB@38_mAd116_1 CB@38_mAd116_2 CB@38_mAd117_1 CB@38_mAd117_2 CB@38_mAd120_1 CB@38_mAd120_2 CB@38_mAd121_1 
+CB@38_mAd121_2 CB@38_mAd122_1 CB@38_mAd122_2 CB@38_mAd123_1 CB@38_mAd123_2 CB@38_mAd124_1 CB@38_mAd124_2 CB@38_mAd125_1 CB@38_mAd125_2 CB@38_mAd126_1 CB@38_mAd126_2 CB@38_mAd127_1 CB@38_mAd127_2 CB@38_mAd130_1 CB@38_mAd130_2 CB@38_mAd131_1 CB@38_mAd131_2 CB@38_mAd132_1 CB@38_mAd132_2 CB@38_mAd133_1 CB@38_mAd133_2 CB@38_mAd134_1 CB@38_mAd134_2 CB@38_mAd135_1 CB@38_mAd135_2 CB@38_mAd136_1 CB@38_mAd136_2 CB@38_mAd137_1 CB@38_mAd137_2 CB@38_mAd140_1 CB@38_mAd140_2 CB@38_mAd141_1 CB@38_mAd141_2 CB@38_mAd142_1 
+CB@38_mAd142_2 CB@38_mAd143_1 CB@38_mAd143_2 CB@38_mAd144_1 CB@38_mAd144_2 CB@38_mAd145_1 CB@38_mAd145_2 CB@38_mAd146_1 CB@38_mAd146_2 CB@38_mAd147_1 CB@38_mAd147_2 CB@38_mAd150_1 CB@38_mAd150_2 CB@38_mAd151_1 CB@38_mAd151_2 CB@38_mAd152_1 CB@38_mAd152_2 CB@38_mAd153_1 CB@38_mAd153_2 CB@38_mAd154_1 CB@38_mAd154_2 CB@38_mAd155_1 CB@38_mAd155_2 CB@38_mAd156_1 CB@38_mAd156_2 CB@38_mAd157_1 CB@38_mAd157_2 CB@38_mAd160_1 CB@38_mAd160_2 CB@38_mAd161_1 CB@38_mAd161_2 CB@38_mAd162_1 CB@38_mAd162_2 CB@38_mAd163_1 
+CB@38_mAd163_2 CB@38_mAd164_1 CB@38_mAd164_2 CB@38_mAd165_1 CB@38_mAd165_2 CB@38_mAd166_1 CB@38_mAd166_2 CB@38_mAd167_1 CB@38_mAd167_2 CB@38_mAd170_1 CB@38_mAd170_2 CB@38_mAd171_1 CB@38_mAd171_2 CB@38_mAd172_1 CB@38_mAd172_2 CB@38_mAd173_1 CB@38_mAd173_2 CB@38_mAd175_1 CB@38_mAd175_2 CB@38_mAd176_1 CB@38_mAd176_2 CB@38_mAd177_1 CB@38_mAd177_2 CB@38_mAd200_1 CB@38_mAd200_2 CB@38_mAd201_1 CB@38_mAd201_2 CB@38_mAd202_1 CB@38_mAd202_2 CB@38_mAd204_1 CB@38_mAd204_2 CB@38_mAd205_1 CB@38_mAd205_2 CB@38_mAd206_1 
+CB@38_mAd206_2 CB@38_mAd207_1 CB@38_mAd207_2 CB@38_mAd210_1 CB@38_mAd210_2 CB@38_mAd211_1 CB@38_mAd211_2 CB@38_mAd212_1 CB@38_mAd212_2 CB@38_mAd213_1 CB@38_mAd213_2 CB@38_mAd214_1 CB@38_mAd214_2 CB@38_mAd215_1 CB@38_mAd215_2 CB@38_mAd216_1 CB@38_mAd216_2 CB@38_mAd217_1 CB@38_mAd217_2 CB@38_mAd220_1 CB@38_mAd220_2 CB@38_mAd221_1 CB@38_mAd221_2 CB@38_mAd222_1 CB@38_mAd222_2 CB@38_mAd223_1 CB@38_mAd223_2 CB@38_mAd224_1 CB@38_mAd224_2 CB@38_mAd225_1 CB@38_mAd225_2 CB@38_mAd226_1 CB@38_mAd226_2 CB@38_mAd227_1 
+CB@38_mAd227_2 CB@38_mAd230_1 CB@38_mAd230_2 CB@38_mAd231_1 CB@38_mAd231_2 CB@38_mAd232_1 CB@38_mAd232_2 CB@38_mAd233_1 CB@38_mAd233_2 CB@38_mAd234_1 CB@38_mAd234_2 CB@38_mAd235_1 CB@38_mAd235_2 CB@38_mAd236_1 CB@38_mAd236_2 CB@38_mAd237_1 CB@38_mAd237_2 CB@38_mAd240_1 CB@38_mAd240_2 CB@38_mAd241_1 CB@38_mAd241_2 CB@38_mAd242_1 CB@38_mAd242_2 CB@38_mAd243_1 CB@38_mAd243_2 CB@38_mAd244_1 CB@38_mAd244_2 CB@38_mAd245_1 CB@38_mAd245_2 CB@38_mAd246_1 CB@38_mAd246_2 CB@38_mAd247_1 CB@38_mAd247_2 CB@38_mAd250_1 
+CB@38_mAd250_2 CB@38_mAd251_1 CB@38_mAd251_2 CB@38_mAd252_1 CB@38_mAd252_2 CB@38_mAd253_1 CB@38_mAd253_2 CB@38_mAd254_1 CB@38_mAd254_2 CB@38_mAd255_1 CB@38_mAd255_2 CB@38_mAd256_1 CB@38_mAd256_2 CB@38_mAd257_1 CB@38_mAd257_2 CB@38_mAd260_1 CB@38_mAd260_2 CB@38_mAd261_1 CB@38_mAd261_2 CB@38_mAd262_1 CB@38_mAd262_2 CB@38_mAd263_1 CB@38_mAd263_2 CB@38_mAd264_1 CB@38_mAd264_2 CB@38_mAd265_1 CB@38_mAd265_2 CB@38_mAd266_1 CB@38_mAd266_2 CB@38_mAd267_1 CB@38_mAd267_2 CB@38_mAd275_1 CB@38_mAd275_2 CB@38_mAd276_1 
+CB@38_mAd276_2 CB@38_mAd277_1 CB@38_mAd277_2 CB@38_mAd300_1 CB@38_mAd300_2 CB@38_mAd310_1 CB@38_mAd310_2 CB@38_mAd311_1 CB@38_mAd311_2 CB@38_mAd317_1 CB@38_mAd317_2 CB@38_mAd320_1 CB@38_mAd320_2 CB@38_mAd321_1 CB@38_mAd321_2 CB@38_mAd322_1 CB@38_mAd322_2 CB@38_mAd323_1 CB@38_mAd323_2 CB@38_mAd324_1 CB@38_mAd324_2 CB@38_mAd325_1 CB@38_mAd325_2 CB@38_mAd326_1 CB@38_mAd326_2 CB@38_mAd327_1 CB@38_mAd327_2 CB@38_mAd330_1 CB@38_mAd330_2 CB@38_mAd331_1 CB@38_mAd331_2 CB@38_mAd332_1 CB@38_mAd332_2 CB@38_mAd333_1 
+CB@38_mAd333_2 CB@38_mAd334_1 CB@38_mAd334_2 CB@38_mAd335_1 CB@38_mAd335_2 CB@38_mAd336_1 CB@38_mAd336_2 CB@38_mAd337_1 CB@38_mAd337_2 CB@38_mAd340_1 CB@38_mAd340_2 CB@38_mAd341_1 CB@38_mAd341_2 CB@38_mAd342_1 CB@38_mAd342_2 CB@38_mAd343_1 CB@38_mAd343_2 CB@38_mAd344_1 CB@38_mAd344_2 CB@38_mAd345_1 CB@38_mAd345_2 CB@38_mAd346_1 CB@38_mAd346_2 CB@38_mAd347_1 CB@38_mAd347_2 CB@38_mAd350_1 CB@38_mAd350_2 CB@38_mAd351_1 CB@38_mAd351_2 CB@38_mAd352_1 CB@38_mAd352_2 CB@38_mAd353_1 CB@38_mAd353_2 CB@38_mAd354_1 
+CB@38_mAd354_2 CB@38_mAd355_1 CB@38_mAd355_2 CB@38_mAd356_1 CB@38_mAd356_2 CB@38_mAd357_1 CB@38_mAd357_2 CB@38_mAd360_1 CB@38_mAd360_2 CB@38_mAd361_1 CB@38_mAd361_2 CB@38_mAd362_1 CB@38_mAd362_2 CB@38_mAd363_1 CB@38_mAd363_2 CB@38_mAd364_1 CB@38_mAd364_2 CB@38_mAd365_1 CB@38_mAd365_2 CB@38_mAd366_1 CB@38_mAd366_2 CB@38_mAd367_1 CB@38_mAd367_2 CB@38_mAd371_1 CB@38_mAd371_2 CB@38_mAd372_1 CB@38_mAd372_2 CB@38_mAd373_1 CB@38_mAd373_2 CB@38_mAd374_1 CB@38_mAd374_2 CB@38_mAd375_1 CB@38_mAd375_2 CB@38_mAd376_1 
+CB@38_mAd376_2 CB@38_mAd377_1 CB@38_mAd377_2 CB@38_mAd400_1 CB@38_mAd400_2 CB@38_mAd401_1 CB@38_mAd401_2 CB@38_mAd402_1 CB@38_mAd402_2 CB@38_mAd403_1 CB@38_mAd403_2 CB@38_mAd404_1 CB@38_mAd404_2 CB@38_mAd405_1 CB@38_mAd405_2 CB@38_mAd406_1 CB@38_mAd406_2 CB@38_mAd407_1 CB@38_mAd407_2 CB@38_mAd410_1 CB@38_mAd410_2 CB@38_mAd411_1 CB@38_mAd411_2 CB@38_mAd412_1 CB@38_mAd412_2 CB@38_mAd413_1 CB@38_mAd413_2 CB@38_mAd414_1 CB@38_mAd414_2 CB@38_mAd415_1 CB@38_mAd415_2 CB@38_mAd416_1 CB@38_mAd416_2 CB@38_mAd417_1 
+CB@38_mAd417_2 CB@38_mAd420_1 CB@38_mAd420_2 CB@38_mAd421_1 CB@38_mAd421_2 CB@38_mAd422_1 CB@38_mAd422_2 CB@38_mAd423_1 CB@38_mAd423_2 CB@38_mAd424_1 CB@38_mAd424_2 CB@38_mAd425_1 CB@38_mAd425_2 CB@38_mAd426_1 CB@38_mAd426_2 CB@38_mAd427_1 CB@38_mAd427_2 CB@38_mAd430_1 CB@38_mAd430_2 CB@38_mAd431_1 CB@38_mAd431_2 CB@38_mAd432_1 CB@38_mAd432_2 CB@38_mAd433_1 CB@38_mAd433_2 CB@38_mAd434_1 CB@38_mAd434_2 CB@38_mAd435_1 CB@38_mAd435_2 CB@38_mAd436_1 CB@38_mAd436_2 CB@38_mAd437_1 CB@38_mAd437_2 CB@38_mAd440_1 
+CB@38_mAd440_2 CB@38_mAd441_1 CB@38_mAd441_2 CB@38_mAd442_1 CB@38_mAd442_2 CB@38_mAd443_1 CB@38_mAd443_2 CB@38_mAd444_1 CB@38_mAd444_2 CB@38_mAd445_1 CB@38_mAd445_2 CB@38_mAd446_1 CB@38_mAd446_2 CB@38_mAd447_1 CB@38_mAd447_2 CB@38_mAd450_1 CB@38_mAd450_2 CB@38_mAd451_1 CB@38_mAd451_2 CB@38_mAd452_1 CB@38_mAd452_2 CB@38_mAd453_1 CB@38_mAd453_2 CB@38_mAd454_1 CB@38_mAd454_2 CB@38_mAd455_1 CB@38_mAd455_2 CB@38_mAd456_1 CB@38_mAd456_2 CB@38_mAd457_1 CB@38_mAd457_2 CB@38_mAd460_1 CB@38_mAd460_2 CB@38_mAd466_1 
+CB@38_mAd466_2 CB@38_mAd467_1 CB@38_mAd467_2 CB@38_mAd500_1 CB@38_mAd500_2 CB@38_mAd501_1 CB@38_mAd501_2 CB@38_mAd502_1 CB@38_mAd502_2 CB@38_mAd508_1 CB@38_mAd508_2 CB@38_mAd509_1 CB@38_mAd509_2 CB@38_mAd512_1 CB@38_mAd512_2 CB@38_mAd513_1 CB@38_mAd513_2 CB@38_mAd514_1 CB@38_mAd514_2 CB@38_mAd515_1 CB@38_mAd515_2 CB@38_mAd516_1 CB@38_mAd516_2 CB@38_mAd517_1 CB@38_mAd517_2 CB@38_mAd520_1 CB@38_mAd520_2 CB@38_mAd521_1 CB@38_mAd521_2 CB@38_mAd522_1 CB@38_mAd522_2 CB@38_mAd523_1 CB@38_mAd523_2 CB@38_mAd524_1 
+CB@38_mAd524_2 CB@38_mAd525_1 CB@38_mAd525_2 CB@38_mAd526_1 CB@38_mAd526_2 CB@38_mAd527_1 CB@38_mAd527_2 CB@38_mAd530_1 CB@38_mAd530_2 CB@38_mAd531_1 CB@38_mAd531_2 CB@38_mAd532_1 CB@38_mAd532_2 CB@38_mAd533_1 CB@38_mAd533_2 CB@38_mAd534_1 CB@38_mAd534_2 CB@38_mAd535_1 CB@38_mAd535_2 CB@38_mAd536_1 CB@38_mAd536_2 CB@38_mAd537_1 CB@38_mAd537_2 CB@38_mAd540_1 CB@38_mAd540_2 CB@38_mAd541_1 CB@38_mAd541_2 CB@38_mAd542_1 CB@38_mAd542_2 CB@38_mAd543_1 CB@38_mAd543_2 CB@38_mAd544_1 CB@38_mAd544_2 CB@38_mAd545_1 
+CB@38_mAd545_2 CB@38_mAd546_1 CB@38_mAd546_2 CB@38_mAd547_1 CB@38_mAd547_2 CB@38_mAd550_1 CB@38_mAd550_2 CB@38_mAd551_1 CB@38_mAd551_2 CB@38_mAd552_1 CB@38_mAd552_2 CB@38_mAd553_1 CB@38_mAd553_2 CB@38_mAd554_1 CB@38_mAd554_2 CB@38_mAd555_1 CB@38_mAd555_2 CB@38_mAd556_1 CB@38_mAd556_2 CB@38_mAd557_1 CB@38_mAd557_2 CB@38_mAd560_1 CB@38_mAd560_2 CB@38_mAd561_1 CB@38_mAd561_2 CB@38_mAd562_1 CB@38_mAd562_2 CB@38_mAd563_1 CB@38_mAd563_2 CB@38_mAd564_1 CB@38_mAd564_2 CB@38_mAd565_1 CB@38_mAd565_2 CB@38_mAd566_1 
+CB@38_mAd566_2 CB@38_mAd567_1 CB@38_mAd567_2 CB@38_mAd570_1 CB@38_mAd570_2 CB@38_mAd571_1 CB@38_mAd571_2 CB@38_mAd572_1 CB@38_mAd572_2 CB@38_mAd573_1 CB@38_mAd573_2 CB@38_mAd575_1 CB@38_mAd575_2 CB@38_mAd576_1 CB@38_mAd576_2 CB@38_mAd577_1 CB@38_mAd577_2 CB@38_mAd600_1 CB@38_mAd600_2 CB@38_mAd601_1 CB@38_mAd601_2 CB@38_mAd602_1 CB@38_mAd602_2 CB@38_mAd604_1 CB@38_mAd604_2 CB@38_mAd605_1 CB@38_mAd605_2 CB@38_mAd606_1 CB@38_mAd606_2 CB@38_mAd607_1 CB@38_mAd607_2 CB@38_mAd610_1 CB@38_mAd610_2 CB@38_mAd611_1 
+CB@38_mAd611_2 CB@38_mAd612_1 CB@38_mAd612_2 CB@38_mAd613_1 CB@38_mAd613_2 CB@38_mAd614_1 CB@38_mAd614_2 CB@38_mAd615_1 CB@38_mAd615_2 CB@38_mAd616_1 CB@38_mAd616_2 CB@38_mAd617_1 CB@38_mAd617_2 CB@38_mAd620_1 CB@38_mAd620_2 CB@38_mAd621_1 CB@38_mAd621_2 CB@38_mAd622_1 CB@38_mAd622_2 CB@38_mAd623_1 CB@38_mAd623_2 CB@38_mAd624_1 CB@38_mAd624_2 CB@38_mAd625_1 CB@38_mAd625_2 CB@38_mAd626_1 CB@38_mAd626_2 CB@38_mAd627_1 CB@38_mAd627_2 CB@38_mAd630_1 CB@38_mAd630_2 CB@38_mAd631_1 CB@38_mAd631_2 CB@38_mAd632_1 
+CB@38_mAd632_2 CB@38_mAd633_1 CB@38_mAd633_2 CB@38_mAd634_1 CB@38_mAd634_2 CB@38_mAd635_1 CB@38_mAd635_2 CB@38_mAd636_1 CB@38_mAd636_2 CB@38_mAd637_1 CB@38_mAd637_2 CB@38_mAd640_1 CB@38_mAd640_2 CB@38_mAd641_1 CB@38_mAd641_2 CB@38_mAd642_1 CB@38_mAd642_2 CB@38_mAd643_1 CB@38_mAd643_2 CB@38_mAd644_1 CB@38_mAd644_2 CB@38_mAd645_1 CB@38_mAd645_2 CB@38_mAd646_1 CB@38_mAd646_2 CB@38_mAd647_1 CB@38_mAd647_2 CB@38_mAd650_1 CB@38_mAd650_2 CB@38_mAd651_1 CB@38_mAd651_2 CB@38_mAd652_1 CB@38_mAd652_2 CB@38_mAd653_1 
+CB@38_mAd653_2 CB@38_mAd654_1 CB@38_mAd654_2 CB@38_mAd655_1 CB@38_mAd655_2 CB@38_mAd656_1 CB@38_mAd656_2 CB@38_mAd657_1 CB@38_mAd657_2 CB@38_mAd660_1 CB@38_mAd660_2 CB@38_mAd661_1 CB@38_mAd661_2 CB@38_mAd662_1 CB@38_mAd662_2 CB@38_mAd663_1 CB@38_mAd663_2 CB@38_mAd664_1 CB@38_mAd664_2 CB@38_mAd665_1 CB@38_mAd665_2 CB@38_mAd666_1 CB@38_mAd666_2 CB@38_mAd667_1 CB@38_mAd667_2 CB@38_mAd675_1 CB@38_mAd675_2 CB@38_mAd676_1 CB@38_mAd676_2 CB@38_mAd677_1 CB@38_mAd677_2 CB@38_mAd700_1 CB@38_mAd700_2 CB@38_mAd710_1 
+CB@38_mAd710_2 CB@38_mAd711_1 CB@38_mAd711_2 CB@38_mAd717_1 CB@38_mAd717_2 CB@38_mAd720_1 CB@38_mAd720_2 CB@38_mAd721_1 CB@38_mAd721_2 CB@38_mAd722_1 CB@38_mAd722_2 CB@38_mAd723_1 CB@38_mAd723_2 CB@38_mAd724_1 CB@38_mAd724_2 CB@38_mAd725_1 CB@38_mAd725_2 CB@38_mAd726_1 CB@38_mAd726_2 CB@38_mAd727_1 CB@38_mAd727_2 CB@38_mAd730_1 CB@38_mAd730_2 CB@38_mAd731_1 CB@38_mAd731_2 CB@38_mAd732_1 CB@38_mAd732_2 CB@38_mAd733_1 CB@38_mAd733_2 CB@38_mAd734_1 CB@38_mAd734_2 CB@38_mAd735_1 CB@38_mAd735_2 CB@38_mAd736_1 
+CB@38_mAd736_2 CB@38_mAd737_1 CB@38_mAd737_2 CB@38_mAd740_1 CB@38_mAd740_2 CB@38_mAd741_1 CB@38_mAd741_2 CB@38_mAd742_1 CB@38_mAd742_2 CB@38_mAd743_1 CB@38_mAd743_2 CB@38_mAd744_1 CB@38_mAd744_2 CB@38_mAd745_1 CB@38_mAd745_2 CB@38_mAd746_1 CB@38_mAd746_2 CB@38_mAd747_1 CB@38_mAd747_2 CB@38_mAd750_1 CB@38_mAd750_2 CB@38_mAd751_1 CB@38_mAd751_2 CB@38_mAd752_1 CB@38_mAd752_2 CB@38_mAd753_1 CB@38_mAd753_2 CB@38_mAd754_1 CB@38_mAd754_2 CB@38_mAd755_1 CB@38_mAd755_2 CB@38_mAd756_1 CB@38_mAd756_2 CB@38_mAd757_1 
+CB@38_mAd757_2 CB@38_mAd760_1 CB@38_mAd760_2 CB@38_mAd761_1 CB@38_mAd761_2 CB@38_mAd762_1 CB@38_mAd762_2 CB@38_mAd763_1 CB@38_mAd763_2 CB@38_mAd764_1 CB@38_mAd764_2 CB@38_mAd765_1 CB@38_mAd765_2 CB@38_mAd766_1 CB@38_mAd766_2 CB@38_mAd767_1 CB@38_mAd767_2 CB@38_mAd771_1 CB@38_mAd771_2 CB@38_mAd772_1 CB@38_mAd772_2 CB@38_mAd773_1 CB@38_mAd773_2 CB@38_mAd774_1 CB@38_mAd774_2 CB@38_mAd775_1 CB@38_mAd775_2 CB@38_mAd776_1 CB@38_mAd776_2 CB@38_mAd777_1 CB@38_mAd777_2 CB@38_X0 CB@38_X1 CB@38_X10 CB@38_X11 
+CB@38_X12 CB@38_X13 CB@38_X2 CB@38_X3 CB@38_X4 CB@38_X5 CB@38_X6 CB@38_X7 CB@38_X8 CB@38_X9 CB@38_Y1 CB@38_Y10 CB@38_Y11 CB@38_Y12 CB@38_Y2 CB@38_Y3 CB@38_Y4 CB@38_Y5 CB@38_Y6 CB@38_Y7 CB@38_Y8 CB@38_Y9 CB@38_Z1 CB@38_Z10 CB@38_Z11 CB@38_Z12 CB@38_Z2 CB@38_Z3 CB@38_Z4 CB@38_Z5 CB@38_Z6 CB@38_Z7 CB@38_Z8 CB@38_Z9 _5400TP094__CB
XCB@39 CB@39_K0 CB@39_K1 CB@39_K10 CB@39_K11 CB@39_K12 CB@39_K13 CB@39_K2 CB@39_K3 CB@39_K4 CB@39_K5 CB@39_K6 CB@39_K7 CB@39_K8 CB@39_K9 CB@39_mAd000_1 CB@39_mAd000_2 CB@39_mAd001_1 CB@39_mAd001_2 CB@39_mAd002_1 CB@39_mAd002_2 CB@39_mAd003_1 CB@39_mAd003_2 CB@39_mAd004_1 CB@39_mAd004_2 CB@39_mAd005_1 CB@39_mAd005_2 CB@39_mAd006_1 CB@39_mAd006_2 CB@39_mAd007_1 CB@39_mAd007_2 CB@39_mAd010_1 CB@39_mAd010_2 CB@39_mAd011_1 CB@39_mAd011_2 CB@39_mAd012_1 CB@39_mAd012_2 CB@39_mAd013_1 CB@39_mAd013_2 CB@39_mAd014_1 
+CB@39_mAd014_2 CB@39_mAd015_1 CB@39_mAd015_2 CB@39_mAd016_1 CB@39_mAd016_2 CB@39_mAd017_1 CB@39_mAd017_2 CB@39_mAd020_1 CB@39_mAd020_2 CB@39_mAd021_1 CB@39_mAd021_2 CB@39_mAd022_1 CB@39_mAd022_2 CB@39_mAd023_1 CB@39_mAd023_2 CB@39_mAd024_1 CB@39_mAd024_2 CB@39_mAd025_1 CB@39_mAd025_2 CB@39_mAd026_1 CB@39_mAd026_2 CB@39_mAd027_1 CB@39_mAd027_2 CB@39_mAd030_1 CB@39_mAd030_2 CB@39_mAd031_1 CB@39_mAd031_2 CB@39_mAd032_1 CB@39_mAd032_2 CB@39_mAd033_1 CB@39_mAd033_2 CB@39_mAd034_1 CB@39_mAd034_2 CB@39_mAd035_1 
+CB@39_mAd035_2 CB@39_mAd036_1 CB@39_mAd036_2 CB@39_mAd037_1 CB@39_mAd037_2 CB@39_mAd040_1 CB@39_mAd040_2 CB@39_mAd041_1 CB@39_mAd041_2 CB@39_mAd042_1 CB@39_mAd042_2 CB@39_mAd043_1 CB@39_mAd043_2 CB@39_mAd044_1 CB@39_mAd044_2 CB@39_mAd045_1 CB@39_mAd045_2 CB@39_mAd046_1 CB@39_mAd046_2 CB@39_mAd047_1 CB@39_mAd047_2 CB@39_mAd050_1 CB@39_mAd050_2 CB@39_mAd051_1 CB@39_mAd051_2 CB@39_mAd052_1 CB@39_mAd052_2 CB@39_mAd053_1 CB@39_mAd053_2 CB@39_mAd054_1 CB@39_mAd054_2 CB@39_mAd055_1 CB@39_mAd055_2 CB@39_mAd056_1 
+CB@39_mAd056_2 CB@39_mAd057_1 CB@39_mAd057_2 CB@39_mAd060_1 CB@39_mAd060_2 CB@39_mAd066_1 CB@39_mAd066_2 CB@39_mAd067_1 CB@39_mAd067_2 CB@39_mAd100_1 CB@39_mAd100_2 CB@39_mAd101_1 CB@39_mAd101_2 CB@39_mAd102_1 CB@39_mAd102_2 CB@39_mAd110_1 CB@39_mAd110_2 CB@39_mAd111_1 CB@39_mAd111_2 CB@39_mAd112_1 CB@39_mAd112_2 CB@39_mAd113_1 CB@39_mAd113_2 CB@39_mAd114_1 CB@39_mAd114_2 CB@39_mAd115_1 CB@39_mAd115_2 CB@39_mAd116_1 CB@39_mAd116_2 CB@39_mAd117_1 CB@39_mAd117_2 CB@39_mAd120_1 CB@39_mAd120_2 CB@39_mAd121_1 
+CB@39_mAd121_2 CB@39_mAd122_1 CB@39_mAd122_2 CB@39_mAd123_1 CB@39_mAd123_2 CB@39_mAd124_1 CB@39_mAd124_2 CB@39_mAd125_1 CB@39_mAd125_2 CB@39_mAd126_1 CB@39_mAd126_2 CB@39_mAd127_1 CB@39_mAd127_2 CB@39_mAd130_1 CB@39_mAd130_2 CB@39_mAd131_1 CB@39_mAd131_2 CB@39_mAd132_1 CB@39_mAd132_2 CB@39_mAd133_1 CB@39_mAd133_2 CB@39_mAd134_1 CB@39_mAd134_2 CB@39_mAd135_1 CB@39_mAd135_2 CB@39_mAd136_1 CB@39_mAd136_2 CB@39_mAd137_1 CB@39_mAd137_2 CB@39_mAd140_1 CB@39_mAd140_2 CB@39_mAd141_1 CB@39_mAd141_2 CB@39_mAd142_1 
+CB@39_mAd142_2 CB@39_mAd143_1 CB@39_mAd143_2 CB@39_mAd144_1 CB@39_mAd144_2 CB@39_mAd145_1 CB@39_mAd145_2 CB@39_mAd146_1 CB@39_mAd146_2 CB@39_mAd147_1 CB@39_mAd147_2 CB@39_mAd150_1 CB@39_mAd150_2 CB@39_mAd151_1 CB@39_mAd151_2 CB@39_mAd152_1 CB@39_mAd152_2 CB@39_mAd153_1 CB@39_mAd153_2 CB@39_mAd154_1 CB@39_mAd154_2 CB@39_mAd155_1 CB@39_mAd155_2 CB@39_mAd156_1 CB@39_mAd156_2 CB@39_mAd157_1 CB@39_mAd157_2 CB@39_mAd160_1 CB@39_mAd160_2 CB@39_mAd161_1 CB@39_mAd161_2 CB@39_mAd162_1 CB@39_mAd162_2 CB@39_mAd163_1 
+CB@39_mAd163_2 CB@39_mAd164_1 CB@39_mAd164_2 CB@39_mAd165_1 CB@39_mAd165_2 CB@39_mAd166_1 CB@39_mAd166_2 CB@39_mAd167_1 CB@39_mAd167_2 CB@39_mAd170_1 CB@39_mAd170_2 CB@39_mAd171_1 CB@39_mAd171_2 CB@39_mAd172_1 CB@39_mAd172_2 CB@39_mAd173_1 CB@39_mAd173_2 CB@39_mAd175_1 CB@39_mAd175_2 CB@39_mAd176_1 CB@39_mAd176_2 CB@39_mAd177_1 CB@39_mAd177_2 CB@39_mAd200_1 CB@39_mAd200_2 CB@39_mAd201_1 CB@39_mAd201_2 CB@39_mAd202_1 CB@39_mAd202_2 CB@39_mAd204_1 CB@39_mAd204_2 CB@39_mAd205_1 CB@39_mAd205_2 CB@39_mAd206_1 
+CB@39_mAd206_2 CB@39_mAd207_1 CB@39_mAd207_2 CB@39_mAd210_1 CB@39_mAd210_2 CB@39_mAd211_1 CB@39_mAd211_2 CB@39_mAd212_1 CB@39_mAd212_2 CB@39_mAd213_1 CB@39_mAd213_2 CB@39_mAd214_1 CB@39_mAd214_2 CB@39_mAd215_1 CB@39_mAd215_2 CB@39_mAd216_1 CB@39_mAd216_2 CB@39_mAd217_1 CB@39_mAd217_2 CB@39_mAd220_1 CB@39_mAd220_2 CB@39_mAd221_1 CB@39_mAd221_2 CB@39_mAd222_1 CB@39_mAd222_2 CB@39_mAd223_1 CB@39_mAd223_2 CB@39_mAd224_1 CB@39_mAd224_2 CB@39_mAd225_1 CB@39_mAd225_2 CB@39_mAd226_1 CB@39_mAd226_2 CB@39_mAd227_1 
+CB@39_mAd227_2 CB@39_mAd230_1 CB@39_mAd230_2 CB@39_mAd231_1 CB@39_mAd231_2 CB@39_mAd232_1 CB@39_mAd232_2 CB@39_mAd233_1 CB@39_mAd233_2 CB@39_mAd234_1 CB@39_mAd234_2 CB@39_mAd235_1 CB@39_mAd235_2 CB@39_mAd236_1 CB@39_mAd236_2 CB@39_mAd237_1 CB@39_mAd237_2 CB@39_mAd240_1 CB@39_mAd240_2 CB@39_mAd241_1 CB@39_mAd241_2 CB@39_mAd242_1 CB@39_mAd242_2 CB@39_mAd243_1 CB@39_mAd243_2 CB@39_mAd244_1 CB@39_mAd244_2 CB@39_mAd245_1 CB@39_mAd245_2 CB@39_mAd246_1 CB@39_mAd246_2 CB@39_mAd247_1 CB@39_mAd247_2 CB@39_mAd250_1 
+CB@39_mAd250_2 CB@39_mAd251_1 CB@39_mAd251_2 CB@39_mAd252_1 CB@39_mAd252_2 CB@39_mAd253_1 CB@39_mAd253_2 CB@39_mAd254_1 CB@39_mAd254_2 CB@39_mAd255_1 CB@39_mAd255_2 CB@39_mAd256_1 CB@39_mAd256_2 CB@39_mAd257_1 CB@39_mAd257_2 CB@39_mAd260_1 CB@39_mAd260_2 CB@39_mAd261_1 CB@39_mAd261_2 CB@39_mAd262_1 CB@39_mAd262_2 CB@39_mAd263_1 CB@39_mAd263_2 CB@39_mAd264_1 CB@39_mAd264_2 CB@39_mAd265_1 CB@39_mAd265_2 CB@39_mAd266_1 CB@39_mAd266_2 CB@39_mAd267_1 CB@39_mAd267_2 CB@39_mAd275_1 CB@39_mAd275_2 CB@39_mAd276_1 
+CB@39_mAd276_2 CB@39_mAd277_1 CB@39_mAd277_2 CB@39_mAd300_1 CB@39_mAd300_2 CB@39_mAd310_1 CB@39_mAd310_2 CB@39_mAd311_1 CB@39_mAd311_2 CB@39_mAd317_1 CB@39_mAd317_2 CB@39_mAd320_1 CB@39_mAd320_2 CB@39_mAd321_1 CB@39_mAd321_2 CB@39_mAd322_1 CB@39_mAd322_2 CB@39_mAd323_1 CB@39_mAd323_2 CB@39_mAd324_1 CB@39_mAd324_2 CB@39_mAd325_1 CB@39_mAd325_2 CB@39_mAd326_1 CB@39_mAd326_2 CB@39_mAd327_1 CB@39_mAd327_2 CB@39_mAd330_1 CB@39_mAd330_2 CB@39_mAd331_1 CB@39_mAd331_2 CB@39_mAd332_1 CB@39_mAd332_2 CB@39_mAd333_1 
+CB@39_mAd333_2 CB@39_mAd334_1 CB@39_mAd334_2 CB@39_mAd335_1 CB@39_mAd335_2 CB@39_mAd336_1 CB@39_mAd336_2 CB@39_mAd337_1 CB@39_mAd337_2 CB@39_mAd340_1 CB@39_mAd340_2 CB@39_mAd341_1 CB@39_mAd341_2 CB@39_mAd342_1 CB@39_mAd342_2 CB@39_mAd343_1 CB@39_mAd343_2 CB@39_mAd344_1 CB@39_mAd344_2 CB@39_mAd345_1 CB@39_mAd345_2 CB@39_mAd346_1 CB@39_mAd346_2 CB@39_mAd347_1 CB@39_mAd347_2 CB@39_mAd350_1 CB@39_mAd350_2 CB@39_mAd351_1 CB@39_mAd351_2 CB@39_mAd352_1 CB@39_mAd352_2 CB@39_mAd353_1 CB@39_mAd353_2 CB@39_mAd354_1 
+CB@39_mAd354_2 CB@39_mAd355_1 CB@39_mAd355_2 CB@39_mAd356_1 CB@39_mAd356_2 CB@39_mAd357_1 CB@39_mAd357_2 CB@39_mAd360_1 CB@39_mAd360_2 CB@39_mAd361_1 CB@39_mAd361_2 CB@39_mAd362_1 CB@39_mAd362_2 CB@39_mAd363_1 CB@39_mAd363_2 CB@39_mAd364_1 CB@39_mAd364_2 CB@39_mAd365_1 CB@39_mAd365_2 CB@39_mAd366_1 CB@39_mAd366_2 CB@39_mAd367_1 CB@39_mAd367_2 CB@39_mAd371_1 CB@39_mAd371_2 CB@39_mAd372_1 CB@39_mAd372_2 CB@39_mAd373_1 CB@39_mAd373_2 CB@39_mAd374_1 CB@39_mAd374_2 CB@39_mAd375_1 CB@39_mAd375_2 CB@39_mAd376_1 
+CB@39_mAd376_2 CB@39_mAd377_1 CB@39_mAd377_2 CB@39_mAd400_1 CB@39_mAd400_2 CB@39_mAd401_1 CB@39_mAd401_2 CB@39_mAd402_1 CB@39_mAd402_2 CB@39_mAd403_1 CB@39_mAd403_2 CB@39_mAd404_1 CB@39_mAd404_2 CB@39_mAd405_1 CB@39_mAd405_2 CB@39_mAd406_1 CB@39_mAd406_2 CB@39_mAd407_1 CB@39_mAd407_2 CB@39_mAd410_1 CB@39_mAd410_2 CB@39_mAd411_1 CB@39_mAd411_2 CB@39_mAd412_1 CB@39_mAd412_2 CB@39_mAd413_1 CB@39_mAd413_2 CB@39_mAd414_1 CB@39_mAd414_2 CB@39_mAd415_1 CB@39_mAd415_2 CB@39_mAd416_1 CB@39_mAd416_2 CB@39_mAd417_1 
+CB@39_mAd417_2 CB@39_mAd420_1 CB@39_mAd420_2 CB@39_mAd421_1 CB@39_mAd421_2 CB@39_mAd422_1 CB@39_mAd422_2 CB@39_mAd423_1 CB@39_mAd423_2 CB@39_mAd424_1 CB@39_mAd424_2 CB@39_mAd425_1 CB@39_mAd425_2 CB@39_mAd426_1 CB@39_mAd426_2 CB@39_mAd427_1 CB@39_mAd427_2 CB@39_mAd430_1 CB@39_mAd430_2 CB@39_mAd431_1 CB@39_mAd431_2 CB@39_mAd432_1 CB@39_mAd432_2 CB@39_mAd433_1 CB@39_mAd433_2 CB@39_mAd434_1 CB@39_mAd434_2 CB@39_mAd435_1 CB@39_mAd435_2 CB@39_mAd436_1 CB@39_mAd436_2 CB@39_mAd437_1 CB@39_mAd437_2 CB@39_mAd440_1 
+CB@39_mAd440_2 CB@39_mAd441_1 CB@39_mAd441_2 CB@39_mAd442_1 CB@39_mAd442_2 CB@39_mAd443_1 CB@39_mAd443_2 CB@39_mAd444_1 CB@39_mAd444_2 CB@39_mAd445_1 CB@39_mAd445_2 CB@39_mAd446_1 CB@39_mAd446_2 CB@39_mAd447_1 CB@39_mAd447_2 CB@39_mAd450_1 CB@39_mAd450_2 CB@39_mAd451_1 CB@39_mAd451_2 CB@39_mAd452_1 CB@39_mAd452_2 CB@39_mAd453_1 CB@39_mAd453_2 CB@39_mAd454_1 CB@39_mAd454_2 CB@39_mAd455_1 CB@39_mAd455_2 CB@39_mAd456_1 CB@39_mAd456_2 CB@39_mAd457_1 CB@39_mAd457_2 CB@39_mAd460_1 CB@39_mAd460_2 CB@39_mAd466_1 
+CB@39_mAd466_2 CB@39_mAd467_1 CB@39_mAd467_2 CB@39_mAd500_1 CB@39_mAd500_2 CB@39_mAd501_1 CB@39_mAd501_2 CB@39_mAd502_1 CB@39_mAd502_2 CB@39_mAd508_1 CB@39_mAd508_2 CB@39_mAd509_1 CB@39_mAd509_2 CB@39_mAd512_1 CB@39_mAd512_2 CB@39_mAd513_1 CB@39_mAd513_2 CB@39_mAd514_1 CB@39_mAd514_2 CB@39_mAd515_1 CB@39_mAd515_2 CB@39_mAd516_1 CB@39_mAd516_2 CB@39_mAd517_1 CB@39_mAd517_2 CB@39_mAd520_1 CB@39_mAd520_2 CB@39_mAd521_1 CB@39_mAd521_2 CB@39_mAd522_1 CB@39_mAd522_2 CB@39_mAd523_1 CB@39_mAd523_2 CB@39_mAd524_1 
+CB@39_mAd524_2 CB@39_mAd525_1 CB@39_mAd525_2 CB@39_mAd526_1 CB@39_mAd526_2 CB@39_mAd527_1 CB@39_mAd527_2 CB@39_mAd530_1 CB@39_mAd530_2 CB@39_mAd531_1 CB@39_mAd531_2 CB@39_mAd532_1 CB@39_mAd532_2 CB@39_mAd533_1 CB@39_mAd533_2 CB@39_mAd534_1 CB@39_mAd534_2 CB@39_mAd535_1 CB@39_mAd535_2 CB@39_mAd536_1 CB@39_mAd536_2 CB@39_mAd537_1 CB@39_mAd537_2 CB@39_mAd540_1 CB@39_mAd540_2 CB@39_mAd541_1 CB@39_mAd541_2 CB@39_mAd542_1 CB@39_mAd542_2 CB@39_mAd543_1 CB@39_mAd543_2 CB@39_mAd544_1 CB@39_mAd544_2 CB@39_mAd545_1 
+CB@39_mAd545_2 CB@39_mAd546_1 CB@39_mAd546_2 CB@39_mAd547_1 CB@39_mAd547_2 CB@39_mAd550_1 CB@39_mAd550_2 CB@39_mAd551_1 CB@39_mAd551_2 CB@39_mAd552_1 CB@39_mAd552_2 CB@39_mAd553_1 CB@39_mAd553_2 CB@39_mAd554_1 CB@39_mAd554_2 CB@39_mAd555_1 CB@39_mAd555_2 CB@39_mAd556_1 CB@39_mAd556_2 CB@39_mAd557_1 CB@39_mAd557_2 CB@39_mAd560_1 CB@39_mAd560_2 CB@39_mAd561_1 CB@39_mAd561_2 CB@39_mAd562_1 CB@39_mAd562_2 CB@39_mAd563_1 CB@39_mAd563_2 CB@39_mAd564_1 CB@39_mAd564_2 CB@39_mAd565_1 CB@39_mAd565_2 CB@39_mAd566_1 
+CB@39_mAd566_2 CB@39_mAd567_1 CB@39_mAd567_2 CB@39_mAd570_1 CB@39_mAd570_2 CB@39_mAd571_1 CB@39_mAd571_2 CB@39_mAd572_1 CB@39_mAd572_2 CB@39_mAd573_1 CB@39_mAd573_2 CB@39_mAd575_1 CB@39_mAd575_2 CB@39_mAd576_1 CB@39_mAd576_2 CB@39_mAd577_1 CB@39_mAd577_2 CB@39_mAd600_1 CB@39_mAd600_2 CB@39_mAd601_1 CB@39_mAd601_2 CB@39_mAd602_1 CB@39_mAd602_2 CB@39_mAd604_1 CB@39_mAd604_2 CB@39_mAd605_1 CB@39_mAd605_2 CB@39_mAd606_1 CB@39_mAd606_2 CB@39_mAd607_1 CB@39_mAd607_2 CB@39_mAd610_1 CB@39_mAd610_2 CB@39_mAd611_1 
+CB@39_mAd611_2 CB@39_mAd612_1 CB@39_mAd612_2 CB@39_mAd613_1 CB@39_mAd613_2 CB@39_mAd614_1 CB@39_mAd614_2 CB@39_mAd615_1 CB@39_mAd615_2 CB@39_mAd616_1 CB@39_mAd616_2 CB@39_mAd617_1 CB@39_mAd617_2 CB@39_mAd620_1 CB@39_mAd620_2 CB@39_mAd621_1 CB@39_mAd621_2 CB@39_mAd622_1 CB@39_mAd622_2 CB@39_mAd623_1 CB@39_mAd623_2 CB@39_mAd624_1 CB@39_mAd624_2 CB@39_mAd625_1 CB@39_mAd625_2 CB@39_mAd626_1 CB@39_mAd626_2 CB@39_mAd627_1 CB@39_mAd627_2 CB@39_mAd630_1 CB@39_mAd630_2 CB@39_mAd631_1 CB@39_mAd631_2 CB@39_mAd632_1 
+CB@39_mAd632_2 CB@39_mAd633_1 CB@39_mAd633_2 CB@39_mAd634_1 CB@39_mAd634_2 CB@39_mAd635_1 CB@39_mAd635_2 CB@39_mAd636_1 CB@39_mAd636_2 CB@39_mAd637_1 CB@39_mAd637_2 CB@39_mAd640_1 CB@39_mAd640_2 CB@39_mAd641_1 CB@39_mAd641_2 CB@39_mAd642_1 CB@39_mAd642_2 CB@39_mAd643_1 CB@39_mAd643_2 CB@39_mAd644_1 CB@39_mAd644_2 CB@39_mAd645_1 CB@39_mAd645_2 CB@39_mAd646_1 CB@39_mAd646_2 CB@39_mAd647_1 CB@39_mAd647_2 CB@39_mAd650_1 CB@39_mAd650_2 CB@39_mAd651_1 CB@39_mAd651_2 CB@39_mAd652_1 CB@39_mAd652_2 CB@39_mAd653_1 
+CB@39_mAd653_2 CB@39_mAd654_1 CB@39_mAd654_2 CB@39_mAd655_1 CB@39_mAd655_2 CB@39_mAd656_1 CB@39_mAd656_2 CB@39_mAd657_1 CB@39_mAd657_2 CB@39_mAd660_1 CB@39_mAd660_2 CB@39_mAd661_1 CB@39_mAd661_2 CB@39_mAd662_1 CB@39_mAd662_2 CB@39_mAd663_1 CB@39_mAd663_2 CB@39_mAd664_1 CB@39_mAd664_2 CB@39_mAd665_1 CB@39_mAd665_2 CB@39_mAd666_1 CB@39_mAd666_2 CB@39_mAd667_1 CB@39_mAd667_2 CB@39_mAd675_1 CB@39_mAd675_2 CB@39_mAd676_1 CB@39_mAd676_2 CB@39_mAd677_1 CB@39_mAd677_2 CB@39_mAd700_1 CB@39_mAd700_2 CB@39_mAd710_1 
+CB@39_mAd710_2 CB@39_mAd711_1 CB@39_mAd711_2 CB@39_mAd717_1 CB@39_mAd717_2 CB@39_mAd720_1 CB@39_mAd720_2 CB@39_mAd721_1 CB@39_mAd721_2 CB@39_mAd722_1 CB@39_mAd722_2 CB@39_mAd723_1 CB@39_mAd723_2 CB@39_mAd724_1 CB@39_mAd724_2 CB@39_mAd725_1 CB@39_mAd725_2 CB@39_mAd726_1 CB@39_mAd726_2 CB@39_mAd727_1 CB@39_mAd727_2 CB@39_mAd730_1 CB@39_mAd730_2 CB@39_mAd731_1 CB@39_mAd731_2 CB@39_mAd732_1 CB@39_mAd732_2 CB@39_mAd733_1 CB@39_mAd733_2 CB@39_mAd734_1 CB@39_mAd734_2 CB@39_mAd735_1 CB@39_mAd735_2 CB@39_mAd736_1 
+CB@39_mAd736_2 CB@39_mAd737_1 CB@39_mAd737_2 CB@39_mAd740_1 CB@39_mAd740_2 CB@39_mAd741_1 CB@39_mAd741_2 CB@39_mAd742_1 CB@39_mAd742_2 CB@39_mAd743_1 CB@39_mAd743_2 CB@39_mAd744_1 CB@39_mAd744_2 CB@39_mAd745_1 CB@39_mAd745_2 CB@39_mAd746_1 CB@39_mAd746_2 CB@39_mAd747_1 CB@39_mAd747_2 CB@39_mAd750_1 CB@39_mAd750_2 CB@39_mAd751_1 CB@39_mAd751_2 CB@39_mAd752_1 CB@39_mAd752_2 CB@39_mAd753_1 CB@39_mAd753_2 CB@39_mAd754_1 CB@39_mAd754_2 CB@39_mAd755_1 CB@39_mAd755_2 CB@39_mAd756_1 CB@39_mAd756_2 CB@39_mAd757_1 
+CB@39_mAd757_2 CB@39_mAd760_1 CB@39_mAd760_2 CB@39_mAd761_1 CB@39_mAd761_2 CB@39_mAd762_1 CB@39_mAd762_2 CB@39_mAd763_1 CB@39_mAd763_2 CB@39_mAd764_1 CB@39_mAd764_2 CB@39_mAd765_1 CB@39_mAd765_2 CB@39_mAd766_1 CB@39_mAd766_2 CB@39_mAd767_1 CB@39_mAd767_2 CB@39_mAd771_1 CB@39_mAd771_2 CB@39_mAd772_1 CB@39_mAd772_2 CB@39_mAd773_1 CB@39_mAd773_2 CB@39_mAd774_1 CB@39_mAd774_2 CB@39_mAd775_1 CB@39_mAd775_2 CB@39_mAd776_1 CB@39_mAd776_2 CB@39_mAd777_1 CB@39_mAd777_2 CB@39_X0 CB@39_X1 CB@39_X10 CB@39_X11 
+CB@39_X12 CB@39_X13 CB@39_X2 CB@39_X3 CB@39_X4 CB@39_X5 CB@39_X6 CB@39_X7 CB@39_X8 CB@39_X9 CB@39_Y1 CB@39_Y10 CB@39_Y11 CB@39_Y12 CB@39_Y2 CB@39_Y3 CB@39_Y4 CB@39_Y5 CB@39_Y6 CB@39_Y7 CB@39_Y8 CB@39_Y9 CB@39_Z1 CB@39_Z10 CB@39_Z11 CB@39_Z12 CB@39_Z2 CB@39_Z3 CB@39_Z4 CB@39_Z5 CB@39_Z6 CB@39_Z7 CB@39_Z8 CB@39_Z9 _5400TP094__CB
Vvsource@1 in1 0 pulse ( 0 2.5 0.1n 0.1n 0.1n 1 2 )
.END
