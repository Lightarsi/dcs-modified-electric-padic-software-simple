*** SPICE deck for cell 123{sch} from library 5400TP094
*** Created on Пн сен 10, 2018 15:16:07
*** Last revised on Пн сен 10, 2018 15:44:42
*** Written on Пн сен 10, 2018 16:17:44 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
.options parhier=local

*** SUBCIRCUIT basic__key FROM CELL basic:key{sch}
.SUBCKT basic__key M1 M2 X Y adr=0
** GLOBAL gnd
Rres@4 gnd M2 100k
*
*
*
*
Xswitch_m@2 X Y M2 switch_man
.SUBCKT switch_man X Y man
S1 X Y man 0 switch1 OFF
.model switch1 sw vt=2.5 vh=1 ron=500 roff=1000G
.ENDS switch_man
******************************************************
Vvsource@0 M1 0 5

* Spice Code nodes in cell cell 'basic:key{sch}'
.param adr = 67
.ENDS basic__key

*** SUBCIRCUIT _5400TP094__CB FROM CELL CB{sch}
.SUBCKT _5400TP094__CB K0 K1 K10 K11 K12 K13 K2 K3 K4 K5 K6 K7 K8 K9 mAd000_1 mAd000_2 mAd001_1 mAd001_2 mAd002_1 mAd002_2 mAd003_1 mAd003_2 mAd004_1 mAd004_2 mAd005_1 mAd005_2 mAd006_1 mAd006_2 mAd007_1 mAd007_2 mAd010_1 mAd010_2 mAd011_1 mAd011_2 mAd012_1 mAd012_2 mAd013_1 mAd013_2 mAd014_1 mAd014_2 mAd015_1 mAd015_2 mAd016_1 mAd016_2 mAd017_1 mAd017_2 mAd020_1 mAd020_2 mAd021_1 mAd021_2 mAd022_1 mAd022_2 mAd023_1 mAd023_2 mAd024_1 mAd024_2 mAd025_1 mAd025_2 mAd026_1 mAd026_2 mAd027_1 mAd027_2 mAd030_1 
+mAd030_2 mAd031_1 mAd031_2 mAd032_1 mAd032_2 mAd033_1 mAd033_2 mAd034_1 mAd034_2 mAd035_1 mAd035_2 mAd036_1 mAd036_2 mAd037_1 mAd037_2 mAd040_1 mAd040_2 mAd041_1 mAd041_2 mAd042_1 mAd042_2 mAd043_1 mAd043_2 mAd044_1 mAd044_2 mAd045_1 mAd045_2 mAd046_1 mAd046_2 mAd047_1 mAd047_2 mAd050_1 mAd050_2 mAd051_1 mAd051_2 mAd052_1 mAd052_2 mAd053_1 mAd053_2 mAd054_1 mAd054_2 mAd055_1 mAd055_2 mAd056_1 mAd056_2 mAd057_1 mAd057_2 mAd060_1 mAd060_2 mAd066_1 mAd066_2 mAd067_1 mAd067_2 mAd100_1 mAd100_2 mAd101_1 
+mAd101_2 mAd102_1 mAd102_2 mAd110_1 mAd110_2 mAd111_1 mAd111_2 mAd112_1 mAd112_2 mAd113_1 mAd113_2 mAd114_1 mAd114_2 mAd115_1 mAd115_2 mAd116_1 mAd116_2 mAd117_1 mAd117_2 mAd120_1 mAd120_2 mAd121_1 mAd121_2 mAd122_1 mAd122_2 mAd123_1 mAd123_2 mAd124_1 mAd124_2 mAd125_1 mAd125_2 mAd126_1 mAd126_2 mAd127_1 mAd127_2 mAd130_1 mAd130_2 mAd131_1 mAd131_2 mAd132_1 mAd132_2 mAd133_1 mAd133_2 mAd134_1 mAd134_2 mAd135_1 mAd135_2 mAd136_1 mAd136_2 mAd137_1 mAd137_2 mAd140_1 mAd140_2 mAd141_1 mAd141_2 mAd142_1 
+mAd142_2 mAd143_1 mAd143_2 mAd144_1 mAd144_2 mAd145_1 mAd145_2 mAd146_1 mAd146_2 mAd147_1 mAd147_2 mAd150_1 mAd150_2 mAd151_1 mAd151_2 mAd152_1 mAd152_2 mAd153_1 mAd153_2 mAd154_1 mAd154_2 mAd155_1 mAd155_2 mAd156_1 mAd156_2 mAd157_1 mAd157_2 mAd160_1 mAd160_2 mAd161_1 mAd161_2 mAd162_1 mAd162_2 mAd163_1 mAd163_2 mAd164_1 mAd164_2 mAd165_1 mAd165_2 mAd166_1 mAd166_2 mAd167_1 mAd167_2 mAd170_1 mAd170_2 mAd171_1 mAd171_2 mAd172_1 mAd172_2 mAd173_1 mAd173_2 mAd175_1 mAd175_2 mAd176_1 mAd176_2 mAd177_1 
+mAd177_2 mAd200_1 mAd200_2 mAd201_1 mAd201_2 mAd202_1 mAd202_2 mAd204_1 mAd204_2 mAd205_1 mAd205_2 mAd206_1 mAd206_2 mAd207_1 mAd207_2 mAd210_1 mAd210_2 mAd211_1 mAd211_2 mAd212_1 mAd212_2 mAd213_1 mAd213_2 mAd214_1 mAd214_2 mAd215_1 mAd215_2 mAd216_1 mAd216_2 mAd217_1 mAd217_2 mAd220_1 mAd220_2 mAd221_1 mAd221_2 mAd222_1 mAd222_2 mAd223_1 mAd223_2 mAd224_1 mAd224_2 mAd225_1 mAd225_2 mAd226_1 mAd226_2 mAd227_1 mAd227_2 mAd230_1 mAd230_2 mAd231_1 mAd231_2 mAd232_1 mAd232_2 mAd233_1 mAd233_2 mAd234_1 
+mAd234_2 mAd235_1 mAd235_2 mAd236_1 mAd236_2 mAd237_1 mAd237_2 mAd240_1 mAd240_2 mAd241_1 mAd241_2 mAd242_1 mAd242_2 mAd243_1 mAd243_2 mAd244_1 mAd244_2 mAd245_1 mAd245_2 mAd246_1 mAd246_2 mAd247_1 mAd247_2 mAd250_1 mAd250_2 mAd251_1 mAd251_2 mAd252_1 mAd252_2 mAd253_1 mAd253_2 mAd254_1 mAd254_2 mAd255_1 mAd255_2 mAd256_1 mAd256_2 mAd257_1 mAd257_2 mAd260_1 mAd260_2 mAd261_1 mAd261_2 mAd262_1 mAd262_2 mAd263_1 mAd263_2 mAd264_1 mAd264_2 mAd265_1 mAd265_2 mAd266_1 mAd266_2 mAd267_1 mAd267_2 mAd275_1 
+mAd275_2 mAd276_1 mAd276_2 mAd277_1 mAd277_2 mAd300_1 mAd300_2 mAd310_1 mAd310_2 mAd311_1 mAd311_2 mAd317_1 mAd317_2 mAd320_1 mAd320_2 mAd321_1 mAd321_2 mAd322_1 mAd322_2 mAd323_1 mAd323_2 mAd324_1 mAd324_2 mAd325_1 mAd325_2 mAd326_1 mAd326_2 mAd327_1 mAd327_2 mAd330_1 mAd330_2 mAd331_1 mAd331_2 mAd332_1 mAd332_2 mAd333_1 mAd333_2 mAd334_1 mAd334_2 mAd335_1 mAd335_2 mAd336_1 mAd336_2 mAd337_1 mAd337_2 mAd340_1 mAd340_2 mAd341_1 mAd341_2 mAd342_1 mAd342_2 mAd343_1 mAd343_2 mAd344_1 mAd344_2 mAd345_1 
+mAd345_2 mAd346_1 mAd346_2 mAd347_1 mAd347_2 mAd350_1 mAd350_2 mAd351_1 mAd351_2 mAd352_1 mAd352_2 mAd353_1 mAd353_2 mAd354_1 mAd354_2 mAd355_1 mAd355_2 mAd356_1 mAd356_2 mAd357_1 mAd357_2 mAd360_1 mAd360_2 mAd361_1 mAd361_2 mAd362_1 mAd362_2 mAd363_1 mAd363_2 mAd364_1 mAd364_2 mAd365_1 mAd365_2 mAd366_1 mAd366_2 mAd367_1 mAd367_2 mAd371_1 mAd371_2 mAd372_1 mAd372_2 mAd373_1 mAd373_2 mAd374_1 mAd374_2 mAd375_1 mAd375_2 mAd376_1 mAd376_2 mAd377_1 mAd377_2 mAd400_1 mAd400_2 mAd401_1 mAd401_2 mAd402_1 
+mAd402_2 mAd403_1 mAd403_2 mAd404_1 mAd404_2 mAd405_1 mAd405_2 mAd406_1 mAd406_2 mAd407_1 mAd407_2 mAd410_1 mAd410_2 mAd411_1 mAd411_2 mAd412_1 mAd412_2 mAd413_1 mAd413_2 mAd414_1 mAd414_2 mAd415_1 mAd415_2 mAd416_1 mAd416_2 mAd417_1 mAd417_2 mAd420_1 mAd420_2 mAd421_1 mAd421_2 mAd422_1 mAd422_2 mAd423_1 mAd423_2 mAd424_1 mAd424_2 mAd425_1 mAd425_2 mAd426_1 mAd426_2 mAd427_1 mAd427_2 mAd430_1 mAd430_2 mAd431_1 mAd431_2 mAd432_1 mAd432_2 mAd433_1 mAd433_2 mAd434_1 mAd434_2 mAd435_1 mAd435_2 mAd436_1 
+mAd436_2 mAd437_1 mAd437_2 mAd440_1 mAd440_2 mAd441_1 mAd441_2 mAd442_1 mAd442_2 mAd443_1 mAd443_2 mAd444_1 mAd444_2 mAd445_1 mAd445_2 mAd446_1 mAd446_2 mAd447_1 mAd447_2 mAd450_1 mAd450_2 mAd451_1 mAd451_2 mAd452_1 mAd452_2 mAd453_1 mAd453_2 mAd454_1 mAd454_2 mAd455_1 mAd455_2 mAd456_1 mAd456_2 mAd457_1 mAd457_2 mAd460_1 mAd460_2 mAd466_1 mAd466_2 mAd467_1 mAd467_2 mAd500_1 mAd500_2 mAd501_1 mAd501_2 mAd502_1 mAd502_2 mAd508_1 mAd508_2 mAd509_1 mAd509_2 mAd512_1 mAd512_2 mAd513_1 mAd513_2 mAd514_1 
+mAd514_2 mAd515_1 mAd515_2 mAd516_1 mAd516_2 mAd517_1 mAd517_2 mAd520_1 mAd520_2 mAd521_1 mAd521_2 mAd522_1 mAd522_2 mAd523_1 mAd523_2 mAd524_1 mAd524_2 mAd525_1 mAd525_2 mAd526_1 mAd526_2 mAd527_1 mAd527_2 mAd530_1 mAd530_2 mAd531_1 mAd531_2 mAd532_1 mAd532_2 mAd533_1 mAd533_2 mAd534_1 mAd534_2 mAd535_1 mAd535_2 mAd536_1 mAd536_2 mAd537_1 mAd537_2 mAd540_1 mAd540_2 mAd541_1 mAd541_2 mAd542_1 mAd542_2 mAd543_1 mAd543_2 mAd544_1 mAd544_2 mAd545_1 mAd545_2 mAd546_1 mAd546_2 mAd547_1 mAd547_2 mAd550_1 
+mAd550_2 mAd551_1 mAd551_2 mAd552_1 mAd552_2 mAd553_1 mAd553_2 mAd554_1 mAd554_2 mAd555_1 mAd555_2 mAd556_1 mAd556_2 mAd557_1 mAd557_2 mAd560_1 mAd560_2 mAd561_1 mAd561_2 mAd562_1 mAd562_2 mAd563_1 mAd563_2 mAd564_1 mAd564_2 mAd565_1 mAd565_2 mAd566_1 mAd566_2 mAd567_1 mAd567_2 mAd570_1 mAd570_2 mAd571_1 mAd571_2 mAd572_1 mAd572_2 mAd573_1 mAd573_2 mAd575_1 mAd575_2 mAd576_1 mAd576_2 mAd577_1 mAd577_2 mAd600_1 mAd600_2 mAd601_1 mAd601_2 mAd602_1 mAd602_2 mAd604_1 mAd604_2 mAd605_1 mAd605_2 mAd606_1 
+mAd606_2 mAd607_1 mAd607_2 mAd610_1 mAd610_2 mAd611_1 mAd611_2 mAd612_1 mAd612_2 mAd613_1 mAd613_2 mAd614_1 mAd614_2 mAd615_1 mAd615_2 mAd616_1 mAd616_2 mAd617_1 mAd617_2 mAd620_1 mAd620_2 mAd621_1 mAd621_2 mAd622_1 mAd622_2 mAd623_1 mAd623_2 mAd624_1 mAd624_2 mAd625_1 mAd625_2 mAd626_1 mAd626_2 mAd627_1 mAd627_2 mAd630_1 mAd630_2 mAd631_1 mAd631_2 mAd632_1 mAd632_2 mAd633_1 mAd633_2 mAd634_1 mAd634_2 mAd635_1 mAd635_2 mAd636_1 mAd636_2 mAd637_1 mAd637_2 mAd640_1 mAd640_2 mAd641_1 mAd641_2 mAd642_1 
+mAd642_2 mAd643_1 mAd643_2 mAd644_1 mAd644_2 mAd645_1 mAd645_2 mAd646_1 mAd646_2 mAd647_1 mAd647_2 mAd650_1 mAd650_2 mAd651_1 mAd651_2 mAd652_1 mAd652_2 mAd653_1 mAd653_2 mAd654_1 mAd654_2 mAd655_1 mAd655_2 mAd656_1 mAd656_2 mAd657_1 mAd657_2 mAd660_1 mAd660_2 mAd661_1 mAd661_2 mAd662_1 mAd662_2 mAd663_1 mAd663_2 mAd664_1 mAd664_2 mAd665_1 mAd665_2 mAd666_1 mAd666_2 mAd667_1 mAd667_2 mAd675_1 mAd675_2 mAd676_1 mAd676_2 mAd677_1 mAd677_2 mAd700_1 mAd700_2 mAd710_1 mAd710_2 mAd711_1 mAd711_2 mAd717_1 
+mAd717_2 mAd720_1 mAd720_2 mAd721_1 mAd721_2 mAd722_1 mAd722_2 mAd723_1 mAd723_2 mAd724_1 mAd724_2 mAd725_1 mAd725_2 mAd726_1 mAd726_2 mAd727_1 mAd727_2 mAd730_1 mAd730_2 mAd731_1 mAd731_2 mAd732_1 mAd732_2 mAd733_1 mAd733_2 mAd734_1 mAd734_2 mAd735_1 mAd735_2 mAd736_1 mAd736_2 mAd737_1 mAd737_2 mAd740_1 mAd740_2 mAd741_1 mAd741_2 mAd742_1 mAd742_2 mAd743_1 mAd743_2 mAd744_1 mAd744_2 mAd745_1 mAd745_2 mAd746_1 mAd746_2 mAd747_1 mAd747_2 mAd750_1 mAd750_2 mAd751_1 mAd751_2 mAd752_1 mAd752_2 mAd753_1 
+mAd753_2 mAd754_1 mAd754_2 mAd755_1 mAd755_2 mAd756_1 mAd756_2 mAd757_1 mAd757_2 mAd760_1 mAd760_2 mAd761_1 mAd761_2 mAd762_1 mAd762_2 mAd763_1 mAd763_2 mAd764_1 mAd764_2 mAd765_1 mAd765_2 mAd766_1 mAd766_2 mAd767_1 mAd767_2 mAd771_1 mAd771_2 mAd772_1 mAd772_2 mAd773_1 mAd773_2 mAd774_1 mAd774_2 mAd775_1 mAd775_2 mAd776_1 mAd776_2 mAd777_1 mAd777_2 X0 X1 X10 X11 X12 X13 X2 X3 X4 X5 X6 X7 X8 X9 Y1 Y10 Y11 Y12 Y2 Y3 Y4 Y5 Y6 Y7 Y8 Y9 Z1 Z10 Z11 Z12 Z2 Z3 Z4 Z5 Z6 Z7 Z8 Z9
** GLOBAL gnd
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
*
Xkey@3 mAd067_1 mAd067_2 K0 X0 basic__key adr=67
Xkey@4 mAd056_1 mAd056_2 X1 Y1 basic__key adr=56
Xkey@5 mAd054_1 mAd054_2 Y1 a2 basic__key adr=54
Xkey@6 mAd046_1 mAd046_2 X1 a1 basic__key adr=46
Xkey@8 mAd044_1 mAd044_2 a1 a2 basic__key adr=44
Xkey@9 mAd055_1 mAd055_2 X1 a2 basic__key adr=55
Xkey@10 mAd045_1 mAd045_2 Y1 a1 basic__key adr=45
Xkey@11 mAd066_1 mAd066_2 Y1 X0 basic__key adr=66
Xkey@12 mAd057_1 mAd057_2 K0 X1 basic__key adr=57
Xkey@13 mAd323_1 mAd323_2 a6 Y12 basic__key adr=323
Xkey@14 mAd321_1 mAd321_2 Y12 Z1 basic__key adr=321
Xkey@15 mAd333_1 mAd333_2 a6 a7 basic__key adr=333
Xkey@16 mAd331_1 mAd331_2 a7 Z1 basic__key adr=331
Xkey@17 mAd322_1 mAd322_2 a6 Z1 basic__key adr=322
Xkey@18 mAd332_1 mAd332_2 Y12 a7 basic__key adr=332
Xkey@19 mAd121_1 mAd121_2 a2 Y6 basic__key adr=121
Xkey@20 mAd160_1 mAd160_2 Y6 a4 basic__key adr=160
Xkey@21 mAd111_1 mAd111_2 a2 a3 basic__key adr=111
Xkey@22 mAd150_1 mAd150_2 a3 a4 basic__key adr=150
Xkey@23 mAd100_1 mAd100_2 a2 a4 basic__key adr=100
Xkey@24 mAd171_1 mAd171_2 Y6 a3 basic__key adr=171
Xkey@25 mAd217_1 mAd217_2 a4 Y7 basic__key adr=217
Xkey@26 mAd256_1 mAd256_2 Y7 a6 basic__key adr=256
Xkey@27 mAd227_1 mAd227_2 a4 a5 basic__key adr=227
Xkey@28 mAd266_1 mAd266_2 a5 a6 basic__key adr=266
Xkey@29 mAd277_1 mAd277_2 a4 a6 basic__key adr=277
Xkey@30 mAd206_1 mAd206_2 Y7 a5 basic__key adr=206
Xkey@31 mAd035_1 mAd035_2 X2 Y2 basic__key adr=35
Xkey@32 mAd033_1 mAd033_2 Y2 b2 basic__key adr=33
Xkey@33 mAd025_1 mAd025_2 X2 b1 basic__key adr=25
Xkey@34 mAd023_1 mAd023_2 b1 b2 basic__key adr=23
Xkey@35 mAd034_1 mAd034_2 X2 b2 basic__key adr=34
Xkey@36 mAd024_1 mAd024_2 Y2 b1 basic__key adr=24
Xkey@37 mAd014_1 mAd014_2 X3 Y3 basic__key adr=14
Xkey@38 mAd012_1 mAd012_2 Y3 c2 basic__key adr=12
Xkey@39 mAd004_1 mAd004_2 X3 c1 basic__key adr=4
Xkey@40 mAd002_1 mAd002_2 c1 c2 basic__key adr=2
Xkey@41 mAd013_1 mAd013_2 X3 c2 basic__key adr=13
Xkey@42 mAd003_1 mAd003_2 Y3 c1 basic__key adr=3
Xkey@43 mAd126_1 mAd126_2 d2 c3 basic__key adr=126
Xkey@44 mAd124_1 mAd124_2 c3 d4 basic__key adr=124
Xkey@45 mAd116_1 mAd116_2 d2 d3 basic__key adr=116
Xkey@46 mAd114_1 mAd114_2 d3 d4 basic__key adr=114
Xkey@47 mAd125_1 mAd125_2 d2 d4 basic__key adr=125
Xkey@48 mAd115_1 mAd115_2 c3 d3 basic__key adr=115
Xkey@49 mAd145_1 mAd145_2 e2 b3 basic__key adr=145
Xkey@50 mAd143_1 mAd143_2 b3 e4 basic__key adr=143
Xkey@51 mAd135_1 mAd135_2 e2 e3 basic__key adr=135
Xkey@52 mAd133_1 mAd133_2 e3 e4 basic__key adr=133
Xkey@53 mAd144_1 mAd144_2 e2 e4 basic__key adr=144
Xkey@54 mAd134_1 mAd134_2 b3 e3 basic__key adr=134
Xkey@55 mAd164_1 mAd164_2 f2 a3 basic__key adr=164
Xkey@56 mAd142_1 mAd142_2 a3 f4 basic__key adr=142
Xkey@57 mAd154_1 mAd154_2 f2 f3 basic__key adr=154
Xkey@58 mAd132_1 mAd132_2 f3 f4 basic__key adr=132
Xkey@59 mAd163_1 mAd163_2 f2 f4 basic__key adr=163
Xkey@60 mAd153_1 mAd153_2 a3 f3 basic__key adr=153
Xkey@61 mAd645_1 mAd645_2 g4 f5 basic__key adr=645
Xkey@62 mAd623_1 mAd623_2 f5 g6 basic__key adr=623
Xkey@63 mAd635_1 mAd635_2 g4 g5 basic__key adr=635
Xkey@64 mAd613_1 mAd613_2 g5 g6 basic__key adr=613
Xkey@65 mAd614_1 mAd614_2 g4 g6 basic__key adr=614
Xkey@66 mAd624_1 mAd624_2 f5 g5 basic__key adr=624
Xkey@67 mAd644_1 mAd644_2 h4 e5 basic__key adr=644
Xkey@68 mAd642_1 mAd642_2 e5 h6 basic__key adr=642
Xkey@69 mAd634_1 mAd634_2 h4 h5 basic__key adr=634
Xkey@70 mAd632_1 mAd632_2 h5 h6 basic__key adr=632
Xkey@71 mAd633_1 mAd633_2 h4 h6 basic__key adr=633
Xkey@72 mAd643_1 mAd643_2 e5 h5 basic__key adr=643
Xkey@73 mAd663_1 mAd663_2 i4 d5 basic__key adr=663
Xkey@74 mAd661_1 mAd661_2 d5 i6 basic__key adr=661
Xkey@75 mAd653_1 mAd653_2 i4 i5 basic__key adr=653
Xkey@76 mAd651_1 mAd651_2 i5 i6 basic__key adr=651
Xkey@77 mAd652_1 mAd652_2 i4 i6 basic__key adr=652
Xkey@78 mAd662_1 mAd662_2 d5 i5 basic__key adr=662
Xkey@79 mAd775_1 mAd775_2 j3 i7 basic__key adr=775
Xkey@80 mAd773_1 mAd773_2 i7 Z10 basic__key adr=773
Xkey@81 mAd765_1 mAd765_2 j3 K10 basic__key adr=765
Xkey@82 mAd763_1 mAd763_2 K10 Z10 basic__key adr=763
Xkey@83 mAd764_1 mAd764_2 j3 Z10 basic__key adr=764
Xkey@84 mAd774_1 mAd774_2 i7 K10 basic__key adr=774
Xkey@85 mAd754_1 mAd754_2 k3 h7 basic__key adr=754
Xkey@86 mAd752_1 mAd752_2 h7 Z11 basic__key adr=752
Xkey@87 mAd744_1 mAd744_2 k3 K11 basic__key adr=744
Xkey@88 mAd742_1 mAd742_2 K11 Z11 basic__key adr=742
Xkey@89 mAd743_1 mAd743_2 k3 Z11 basic__key adr=743
Xkey@90 mAd753_1 mAd753_2 h7 K11 basic__key adr=753
Xkey@91 mAd733_1 mAd733_2 l3 g7 basic__key adr=733
Xkey@92 mAd731_1 mAd731_2 g7 Z12 basic__key adr=731
Xkey@93 mAd723_1 mAd723_2 l3 K12 basic__key adr=723
Xkey@94 mAd721_1 mAd721_2 K12 Z12 basic__key adr=721
Xkey@95 mAd722_1 mAd722_2 l3 Z12 basic__key adr=722
Xkey@96 mAd732_1 mAd732_2 g7 K12 basic__key adr=732
Xkey@97 mAd037_1 mAd037_2 K0 X2 basic__key adr=37
Xkey@98 mAd017_1 mAd017_2 K0 X3 basic__key adr=17
Xkey@99 mAd007_1 mAd007_2 K0 X4 basic__key adr=7
Xkey@100 mAd027_1 mAd027_2 K0 X5 basic__key adr=27
Xkey@101 mAd047_1 mAd047_2 K0 X6 basic__key adr=47
Xkey@102 mAd447_1 mAd447_2 K0 X7 basic__key adr=447
Xkey@103 mAd427_1 mAd427_2 K0 X8 basic__key adr=427
Xkey@104 mAd407_1 mAd407_2 K0 X9 basic__key adr=407
Xkey@105 mAd417_1 mAd417_2 K0 X10 basic__key adr=417
Xkey@106 mAd437_1 mAd437_2 K0 X11 basic__key adr=437
Xkey@107 mAd457_1 mAd457_2 K0 X12 basic__key adr=457
Xkey@108 mAd467_1 mAd467_2 K0 X13 basic__key adr=467
Xkey@109 mAd446_1 mAd446_2 X12 g1 basic__key adr=446
Xkey@110 mAd444_1 mAd444_2 g1 l1 basic__key adr=444
Xkey@111 mAd456_1 mAd456_2 X12 K1 basic__key adr=456
Xkey@112 mAd454_1 mAd454_2 K1 l1 basic__key adr=454
Xkey@113 mAd455_1 mAd455_2 X12 l1 basic__key adr=455
Xkey@114 mAd445_1 mAd445_2 g1 K1 basic__key adr=445
Xkey@115 mAd425_1 mAd425_2 X11 h1 basic__key adr=425
Xkey@116 mAd423_1 mAd423_2 h1 k1 basic__key adr=423
Xkey@117 mAd435_1 mAd435_2 X11 K2 basic__key adr=435
Xkey@118 mAd433_1 mAd433_2 K2 k1 basic__key adr=433
Xkey@119 mAd434_1 mAd434_2 X11 k1 basic__key adr=434
Xkey@120 mAd424_1 mAd424_2 h1 K2 basic__key adr=424
Xkey@121 mAd404_1 mAd404_2 X10 i1 basic__key adr=404
Xkey@122 mAd402_1 mAd402_2 i1 j1 basic__key adr=402
Xkey@123 mAd414_1 mAd414_2 X10 K3 basic__key adr=414
Xkey@124 mAd412_1 mAd412_2 K3 j1 basic__key adr=412
Xkey@125 mAd413_1 mAd413_2 X10 j1 basic__key adr=413
Xkey@126 mAd403_1 mAd403_2 i1 K3 basic__key adr=403
Xkey@127 mAd516_1 mAd516_2 i2 d3 basic__key adr=516
Xkey@128 mAd514_1 mAd514_2 d3 i4 basic__key adr=514
Xkey@129 mAd526_1 mAd526_2 i2 i3 basic__key adr=526
Xkey@130 mAd524_1 mAd524_2 i3 i4 basic__key adr=524
Xkey@131 mAd525_1 mAd525_2 i2 i4 basic__key adr=525
Xkey@132 mAd515_1 mAd515_2 d3 i3 basic__key adr=515
Xkey@133 mAd535_1 mAd535_2 h2 e3 basic__key adr=535
Xkey@134 mAd533_1 mAd533_2 e3 h4 basic__key adr=533
Xkey@135 mAd545_1 mAd545_2 h2 h3 basic__key adr=545
Xkey@136 mAd543_1 mAd543_2 h3 h4 basic__key adr=543
Xkey@137 mAd544_1 mAd544_2 h2 h4 basic__key adr=544
Xkey@138 mAd534_1 mAd534_2 e3 h3 basic__key adr=534
Xkey@139 mAd554_1 mAd554_2 g2 f3 basic__key adr=554
Xkey@140 mAd532_1 mAd532_2 f3 g4 basic__key adr=532
Xkey@141 mAd564_1 mAd564_2 g2 g3 basic__key adr=564
Xkey@142 mAd542_1 mAd542_2 g3 g4 basic__key adr=542
Xkey@143 mAd563_1 mAd563_2 g2 g4 basic__key adr=563
Xkey@144 mAd553_1 mAd553_2 f3 g3 basic__key adr=553
Xkey@145 mAd235_1 mAd235_2 f4 a5 basic__key adr=235
Xkey@146 mAd213_1 mAd213_2 a5 f6 basic__key adr=213
Xkey@147 mAd245_1 mAd245_2 f4 f5 basic__key adr=245
Xkey@148 mAd223_1 mAd223_2 f5 f6 basic__key adr=223
Xkey@149 mAd214_1 mAd214_2 f4 f6 basic__key adr=214
Xkey@150 mAd224_1 mAd224_2 a5 f5 basic__key adr=224
Xkey@151 mAd234_1 mAd234_2 e4 b5 basic__key adr=234
Xkey@152 mAd232_1 mAd232_2 b5 e6 basic__key adr=232
Xkey@153 mAd244_1 mAd244_2 e4 e5 basic__key adr=244
Xkey@154 mAd242_1 mAd242_2 e5 e6 basic__key adr=242
Xkey@155 mAd233_1 mAd233_2 e4 e6 basic__key adr=233
Xkey@156 mAd243_1 mAd243_2 b5 e5 basic__key adr=243
Xkey@157 mAd253_1 mAd253_2 d4 c5 basic__key adr=253
Xkey@158 mAd251_1 mAd251_2 c5 d6 basic__key adr=251
Xkey@159 mAd263_1 mAd263_2 d4 d5 basic__key adr=263
Xkey@160 mAd261_1 mAd261_2 d5 d6 basic__key adr=261
Xkey@161 mAd252_1 mAd252_2 d4 d6 basic__key adr=252
Xkey@162 mAd262_1 mAd262_2 c5 d5 basic__key adr=262
Xkey@163 mAd365_1 mAd365_2 c6 Y10 basic__key adr=365
Xkey@164 mAd363_1 mAd363_2 Y10 Z3 basic__key adr=363
Xkey@165 mAd375_1 mAd375_2 c6 c7 basic__key adr=375
Xkey@166 mAd373_1 mAd373_2 c7 Z3 basic__key adr=373
Xkey@167 mAd364_1 mAd364_2 c6 Z3 basic__key adr=364
Xkey@168 mAd374_1 mAd374_2 Y10 c7 basic__key adr=374
Xkey@169 mAd344_1 mAd344_2 b6 Y11 basic__key adr=344
Xkey@170 mAd342_1 mAd342_2 Y11 Z2 basic__key adr=342
Xkey@171 mAd354_1 mAd354_2 b6 b7 basic__key adr=354
Xkey@172 mAd352_1 mAd352_2 b7 Z2 basic__key adr=352
Xkey@173 mAd343_1 mAd343_2 b6 Z2 basic__key adr=343
Xkey@174 mAd353_1 mAd353_2 Y11 b7 basic__key adr=353
Xkey@175 mAd122_1 mAd122_2 b2 Y5 basic__key adr=122
Xkey@176 mAd161_1 mAd161_2 Y5 b4 basic__key adr=161
Xkey@177 mAd112_1 mAd112_2 b2 b3 basic__key adr=112
Xkey@178 mAd151_1 mAd151_2 b3 b4 basic__key adr=151
Xkey@179 mAd101_1 mAd101_2 b2 b4 basic__key adr=101
Xkey@180 mAd172_1 mAd172_2 Y5 b3 basic__key adr=172
Xkey@181 mAd123_1 mAd123_2 c2 Y4 basic__key adr=123
Xkey@182 mAd162_1 mAd162_2 Y4 c4 basic__key adr=162
Xkey@183 mAd113_1 mAd113_2 c2 c3 basic__key adr=113
Xkey@184 mAd152_1 mAd152_2 c3 c4 basic__key adr=152
Xkey@185 mAd102_1 mAd102_2 c2 c4 basic__key adr=102
Xkey@186 mAd173_1 mAd173_2 Y4 c3 basic__key adr=173
Xkey@187 mAd011_1 mAd011_2 X4 c1 basic__key adr=11
Xkey@188 mAd127_1 mAd127_2 c1 d2 basic__key adr=127
Xkey@189 mAd001_1 mAd001_2 X4 d1 basic__key adr=1
Xkey@190 mAd117_1 mAd117_2 d1 d2 basic__key adr=117
Xkey@191 mAd010_1 mAd010_2 X4 d2 basic__key adr=10
Xkey@192 mAd000_1 mAd000_2 c1 d1 basic__key adr=0
Xkey@193 mAd032_1 mAd032_2 X5 b1 basic__key adr=32
Xkey@194 mAd030_1 mAd030_2 b1 e2 basic__key adr=30
Xkey@195 mAd022_1 mAd022_2 X5 e1 basic__key adr=22
Xkey@196 mAd020_1 mAd020_2 e1 e2 basic__key adr=20
Xkey@197 mAd031_1 mAd031_2 X5 e2 basic__key adr=31
Xkey@198 mAd021_1 mAd021_2 b1 e1 basic__key adr=21
Xkey@199 mAd053_1 mAd053_2 X6 a1 basic__key adr=53
Xkey@200 mAd051_1 mAd051_2 a1 f2 basic__key adr=51
Xkey@201 mAd043_1 mAd043_2 X6 f1 basic__key adr=43
Xkey@202 mAd041_1 mAd041_2 f1 f2 basic__key adr=41
Xkey@203 mAd052_1 mAd052_2 X6 f2 basic__key adr=52
Xkey@204 mAd042_1 mAd042_2 a1 f1 basic__key adr=42
Xkey@205 mAd443_1 mAd443_2 X7 f1 basic__key adr=443
Xkey@206 mAd441_1 mAd441_2 f1 g2 basic__key adr=441
Xkey@207 mAd453_1 mAd453_2 X7 g1 basic__key adr=453
Xkey@208 mAd451_1 mAd451_2 g1 g2 basic__key adr=451
Xkey@209 mAd452_1 mAd452_2 X7 g2 basic__key adr=452
Xkey@210 mAd442_1 mAd442_2 f1 g1 basic__key adr=442
Xkey@211 mAd422_1 mAd422_2 X8 e1 basic__key adr=422
Xkey@212 mAd420_1 mAd420_2 e1 h2 basic__key adr=420
Xkey@213 mAd432_1 mAd432_2 X8 h1 basic__key adr=432
Xkey@214 mAd430_1 mAd430_2 h1 h2 basic__key adr=430
Xkey@215 mAd431_1 mAd431_2 X8 h2 basic__key adr=431
Xkey@216 mAd421_1 mAd421_2 e1 h1 basic__key adr=421
Xkey@217 mAd401_1 mAd401_2 X9 d1 basic__key adr=401
Xkey@218 mAd517_1 mAd517_2 d1 i2 basic__key adr=517
Xkey@219 mAd411_1 mAd411_2 X9 i1 basic__key adr=411
Xkey@220 mAd527_1 mAd527_2 i1 i2 basic__key adr=527
Xkey@221 mAd410_1 mAd410_2 X9 i2 basic__key adr=410
Xkey@222 mAd400_1 mAd400_2 d1 i1 basic__key adr=400
Xkey@223 mAd513_1 mAd513_2 j1 i3 basic__key adr=513
Xkey@224 mAd552_1 mAd552_2 i3 j2 basic__key adr=552
Xkey@225 mAd523_1 mAd523_2 j1 K4 basic__key adr=523
Xkey@226 mAd562_1 mAd562_2 K4 j2 basic__key adr=562
Xkey@227 mAd502_1 mAd502_2 j1 j2 basic__key adr=502
Xkey@228 mAd573_1 mAd573_2 i3 K4 basic__key adr=573
Xkey@229 mAd512_1 mAd512_2 k1 h3 basic__key adr=512
Xkey@230 mAd551_1 mAd551_2 h3 k2 basic__key adr=551
Xkey@231 mAd522_1 mAd522_2 k1 K5 basic__key adr=522
Xkey@232 mAd561_1 mAd561_2 K5 k2 basic__key adr=561
Xkey@233 mAd501_1 mAd501_2 k1 k2 basic__key adr=501
Xkey@234 mAd572_1 mAd572_2 h3 K5 basic__key adr=572
Xkey@235 mAd509_1 mAd509_2 l1 g3 basic__key adr=509
Xkey@236 mAd550_1 mAd550_2 g3 l2 basic__key adr=550
Xkey@237 mAd521_1 mAd521_2 l1 K6 basic__key adr=521
Xkey@238 mAd560_1 mAd560_2 K6 l2 basic__key adr=560
Xkey@239 mAd500_1 mAd500_2 l1 l2 basic__key adr=500
Xkey@240 mAd571_1 mAd571_2 g3 K6 basic__key adr=571
Xkey@241 mAd627_1 mAd627_2 l2 g5 basic__key adr=627
Xkey@242 mAd666_1 mAd666_2 g5 l3 basic__key adr=666
Xkey@243 mAd617_1 mAd617_2 l2 K7 basic__key adr=617
Xkey@244 mAd656_1 mAd656_2 K7 l3 basic__key adr=656
Xkey@245 mAd677_1 mAd677_2 l2 l3 basic__key adr=677
Xkey@246 mAd606_1 mAd606_2 g5 K7 basic__key adr=606
Xkey@247 mAd626_1 mAd626_2 k2 h5 basic__key adr=626
Xkey@248 mAd665_1 mAd665_2 h5 k3 basic__key adr=665
Xkey@249 mAd616_1 mAd616_2 k2 K8 basic__key adr=616
Xkey@250 mAd655_1 mAd655_2 K8 k3 basic__key adr=655
Xkey@251 mAd676_1 mAd676_2 k2 k3 basic__key adr=676
Xkey@252 mAd605_1 mAd605_2 h5 K8 basic__key adr=605
Xkey@253 mAd625_1 mAd625_2 j2 i5 basic__key adr=625
Xkey@254 mAd664_1 mAd664_2 i5 j3 basic__key adr=664
Xkey@255 mAd615_1 mAd615_2 j2 K9 basic__key adr=615
Xkey@256 mAd654_1 mAd654_2 K9 j3 basic__key adr=654
Xkey@257 mAd675_1 mAd675_2 j2 j3 basic__key adr=675
Xkey@258 mAd604_1 mAd604_2 i5 K9 basic__key adr=604
Xkey@259 mAd660_1 mAd660_2 i6 d7 basic__key adr=660
Xkey@260 mAd776_1 mAd776_2 d7 Z9 basic__key adr=776
Xkey@261 mAd650_1 mAd650_2 i6 i7 basic__key adr=650
Xkey@262 mAd766_1 mAd766_2 i7 Z9 basic__key adr=766
Xkey@263 mAd767_1 mAd767_2 i6 Z9 basic__key adr=767
Xkey@264 mAd777_1 mAd777_2 d7 i7 basic__key adr=777
Xkey@265 mAd757_1 mAd757_2 h6 e7 basic__key adr=757
Xkey@266 mAd755_1 mAd755_2 e7 Z8 basic__key adr=755
Xkey@267 mAd747_1 mAd747_2 h6 h7 basic__key adr=747
Xkey@268 mAd745_1 mAd745_2 h7 Z8 basic__key adr=745
Xkey@269 mAd746_1 mAd746_2 h6 Z8 basic__key adr=746
Xkey@270 mAd756_1 mAd756_2 e7 h7 basic__key adr=756
Xkey@271 mAd736_1 mAd736_2 g6 f7 basic__key adr=736
Xkey@272 mAd734_1 mAd734_2 f7 Z7 basic__key adr=734
Xkey@273 mAd726_1 mAd726_2 g6 g7 basic__key adr=726
Xkey@274 mAd724_1 mAd724_2 g7 Z7 basic__key adr=724
Xkey@275 mAd725_1 mAd725_2 g6 Z7 basic__key adr=725
Xkey@276 mAd735_1 mAd735_2 f7 g7 basic__key adr=735
Xkey@277 mAd326_1 mAd326_2 f6 a7 basic__key adr=326
Xkey@278 mAd324_1 mAd324_2 a7 Z6 basic__key adr=324
Xkey@279 mAd336_1 mAd336_2 f6 f7 basic__key adr=336
Xkey@280 mAd334_1 mAd334_2 f7 Z6 basic__key adr=334
Xkey@281 mAd325_1 mAd325_2 f6 Z6 basic__key adr=325
Xkey@282 mAd335_1 mAd335_2 a7 f7 basic__key adr=335
Xkey@283 mAd347_1 mAd347_2 e6 b7 basic__key adr=347
Xkey@284 mAd345_1 mAd345_2 b7 Z5 basic__key adr=345
Xkey@285 mAd357_1 mAd357_2 e6 e7 basic__key adr=357
Xkey@286 mAd355_1 mAd355_2 e7 Z5 basic__key adr=355
Xkey@287 mAd346_1 mAd346_2 e6 Z5 basic__key adr=346
Xkey@288 mAd356_1 mAd356_2 b7 e7 basic__key adr=356
Xkey@289 mAd250_1 mAd250_2 d6 c7 basic__key adr=250
Xkey@290 mAd366_1 mAd366_2 c7 Z4 basic__key adr=366
Xkey@291 mAd260_1 mAd260_2 d6 d7 basic__key adr=260
Xkey@292 mAd376_1 mAd376_2 d7 Z4 basic__key adr=376
Xkey@293 mAd367_1 mAd367_2 d6 Z4 basic__key adr=367
Xkey@294 mAd377_1 mAd377_2 c7 d7 basic__key adr=377
Xkey@295 mAd215_1 mAd215_2 c4 Y9 basic__key adr=215
Xkey@296 mAd254_1 mAd254_2 Y9 c6 basic__key adr=254
Xkey@297 mAd225_1 mAd225_2 c4 c5 basic__key adr=225
Xkey@298 mAd264_1 mAd264_2 c5 c6 basic__key adr=264
Xkey@299 mAd275_1 mAd275_2 c4 c6 basic__key adr=275
Xkey@300 mAd204_1 mAd204_2 Y9 c5 basic__key adr=204
Xkey@301 mAd216_1 mAd216_2 b4 Y8 basic__key adr=216
Xkey@302 mAd255_1 mAd255_2 Y8 b6 basic__key adr=255
Xkey@303 mAd226_1 mAd226_2 b4 b5 basic__key adr=226
Xkey@304 mAd265_1 mAd265_2 b5 b6 basic__key adr=265
Xkey@305 mAd276_1 mAd276_2 b4 b6 basic__key adr=276
Xkey@306 mAd205_1 mAd205_2 Y8 b5 basic__key adr=205
Xkey@307 mAd060_1 mAd060_2 Y2 X0 basic__key adr=60
Xkey@308 mAd177_1 mAd177_2 Y3 X0 basic__key adr=177
Xkey@309 mAd176_1 mAd176_2 Y4 X0 basic__key adr=176
Xkey@310 mAd175_1 mAd175_2 Y5 X0 basic__key adr=175
Xkey@311 mAd170_1 mAd170_2 Y6 X0 basic__key adr=170
Xkey@312 mAd207_1 mAd207_2 Y7 X0 basic__key adr=207
Xkey@313 mAd202_1 mAd202_2 Y8 X0 basic__key adr=202
Xkey@314 mAd201_1 mAd201_2 Y9 X0 basic__key adr=201
Xkey@315 mAd200_1 mAd200_2 Y10 X0 basic__key adr=200
Xkey@316 mAd317_1 mAd317_2 Y11 X0 basic__key adr=317
Xkey@317 mAd311_1 mAd311_2 Y12 X0 basic__key adr=311
Xkey@318 mAd300_1 mAd300_2 K13 X0 basic__key adr=300
Xkey@319 mAd050_1 mAd050_2 Y2 a2 basic__key adr=50
Xkey@320 mAd167_1 mAd167_2 Y3 a2 basic__key adr=167
Xkey@321 mAd166_1 mAd166_2 Y4 a2 basic__key adr=166
Xkey@322 mAd165_1 mAd165_2 Y5 a2 basic__key adr=165
Xkey@323 mAd212_1 mAd212_2 Y8 a6 basic__key adr=212
Xkey@324 mAd211_1 mAd211_2 Y9 a6 basic__key adr=211
Xkey@325 mAd210_1 mAd210_2 Y10 a6 basic__key adr=210
Xkey@326 mAd327_1 mAd327_2 Y11 a6 basic__key adr=327
Xkey@327 mAd310_1 mAd310_2 K13 Z1 basic__key adr=310
Xkey@328 mAd036_1 mAd036_2 a1 X2 basic__key adr=36
Xkey@329 mAd147_1 mAd147_2 Y3 b2 basic__key adr=147
Xkey@330 mAd146_1 mAd146_2 Y4 b2 basic__key adr=146
Xkey@331 mAd140_1 mAd140_2 a3 b4 basic__key adr=140
Xkey@332 mAd237_1 mAd237_2 a5 b4 basic__key adr=237
Xkey@333 mAd231_1 mAd231_2 Y9 b6 basic__key adr=231
Xkey@334 mAd230_1 mAd230_2 Y10 b6 basic__key adr=230
Xkey@335 mAd341_1 mAd341_2 a7 Z2 basic__key adr=341
Xkey@336 mAd330_1 mAd330_2 K13 Z2 basic__key adr=330
Xkey@337 mAd016_1 mAd016_2 a1 X3 basic__key adr=16
Xkey@338 mAd015_1 mAd015_2 b1 X3 basic__key adr=15
Xkey@339 mAd141_1 mAd141_2 b3 c4 basic__key adr=141
Xkey@340 mAd120_1 mAd120_2 a3 c4 basic__key adr=120
Xkey@341 mAd257_1 mAd257_2 a5 c4 basic__key adr=257
Xkey@342 mAd236_1 mAd236_2 b5 c4 basic__key adr=236
Xkey@343 mAd362_1 mAd362_2 b7 Z3 basic__key adr=362
Xkey@344 mAd361_1 mAd361_2 a7 Z3 basic__key adr=361
Xkey@345 mAd350_1 mAd350_2 K13 Z3 basic__key adr=350
Xkey@346 mAd360_1 mAd360_2 K13 Z4 basic__key adr=360
Xkey@347 mAd371_1 mAd371_2 a7 Z4 basic__key adr=371
Xkey@348 mAd372_1 mAd372_2 b7 Z4 basic__key adr=372
Xkey@349 mAd246_1 mAd246_2 b5 d4 basic__key adr=246
Xkey@350 mAd267_1 mAd267_2 a5 d4 basic__key adr=267
Xkey@351 mAd110_1 mAd110_2 a3 d4 basic__key adr=110
Xkey@352 mAd131_1 mAd131_2 b3 d4 basic__key adr=131
Xkey@353 mAd005_1 mAd005_2 b1 X4 basic__key adr=5
Xkey@354 mAd006_1 mAd006_2 a1 X4 basic__key adr=6
Xkey@355 mAd026_1 mAd026_2 a1 X5 basic__key adr=26
Xkey@356 mAd137_1 mAd137_2 d1 e2 basic__key adr=137
Xkey@357 mAd136_1 mAd136_2 d3 e2 basic__key adr=136
Xkey@358 mAd130_1 mAd130_2 a3 e4 basic__key adr=130
Xkey@359 mAd247_1 mAd247_2 a5 e4 basic__key adr=247
Xkey@360 mAd241_1 mAd241_2 d5 e6 basic__key adr=241
Xkey@361 mAd240_1 mAd240_2 d7 e6 basic__key adr=240
Xkey@362 mAd351_1 mAd351_2 a7 Z5 basic__key adr=351
Xkey@363 mAd340_1 mAd340_2 K13 Z5 basic__key adr=340
Xkey@364 mAd320_1 mAd320_2 K13 Z6 basic__key adr=320
Xkey@365 mAd337_1 mAd337_2 e7 f6 basic__key adr=337
Xkey@366 mAd220_1 mAd220_2 d7 f6 basic__key adr=220
Xkey@367 mAd221_1 mAd221_2 d5 f6 basic__key adr=221
Xkey@368 mAd222_1 mAd222_2 e5 f6 basic__key adr=222
Xkey@369 mAd155_1 mAd155_2 e3 f2 basic__key adr=155
Xkey@370 mAd156_1 mAd156_2 d3 f2 basic__key adr=156
Xkey@371 mAd157_1 mAd157_2 d1 f2 basic__key adr=157
Xkey@372 mAd040_1 mAd040_2 e1 f2 basic__key adr=40
Xkey@373 mAd440_1 mAd440_2 e1 g2 basic__key adr=440
Xkey@374 mAd557_1 mAd557_2 d1 g2 basic__key adr=557
Xkey@375 mAd556_1 mAd556_2 d3 g2 basic__key adr=556
Xkey@376 mAd555_1 mAd555_2 e3 g2 basic__key adr=555
Xkey@377 mAd622_1 mAd622_2 e5 g6 basic__key adr=622
Xkey@378 mAd621_1 mAd621_2 d5 g6 basic__key adr=621
Xkey@379 mAd620_1 mAd620_2 d7 g6 basic__key adr=620
Xkey@380 mAd737_1 mAd737_2 e7 g6 basic__key adr=737
Xkey@381 mAd720_1 mAd720_2 K13 Z7 basic__key adr=720
Xkey@382 mAd426_1 mAd426_2 g1 X8 basic__key adr=426
Xkey@383 mAd537_1 mAd537_2 d1 h2 basic__key adr=537
Xkey@384 mAd536_1 mAd536_2 d3 h2 basic__key adr=536
Xkey@385 mAd530_1 mAd530_2 g3 h4 basic__key adr=530
Xkey@386 mAd647_1 mAd647_2 g5 h4 basic__key adr=647
Xkey@387 mAd641_1 mAd641_2 d5 h6 basic__key adr=641
Xkey@388 mAd640_1 mAd640_2 d7 h6 basic__key adr=640
Xkey@389 mAd751_1 mAd751_2 g7 Z8 basic__key adr=751
Xkey@390 mAd740_1 mAd740_2 K13 Z8 basic__key adr=740
Xkey@391 mAd406_1 mAd406_2 g1 X9 basic__key adr=406
Xkey@392 mAd405_1 mAd405_2 h1 X9 basic__key adr=405
Xkey@393 mAd531_1 mAd531_2 h3 i4 basic__key adr=531
Xkey@394 mAd508_1 mAd508_2 g3 i4 basic__key adr=508
Xkey@395 mAd667_1 mAd667_2 g5 i4 basic__key adr=667
Xkey@396 mAd646_1 mAd646_2 h5 i4 basic__key adr=646
Xkey@397 mAd772_1 mAd772_2 h7 Z9 basic__key adr=772
Xkey@398 mAd771_1 mAd771_2 g7 Z9 basic__key adr=771
Xkey@399 mAd760_1 mAd760_2 K13 Z9 basic__key adr=760
Xkey@400 mAd416_1 mAd416_2 g1 X10 basic__key adr=416
Xkey@401 mAd415_1 mAd415_2 h1 X10 basic__key adr=415
Xkey@402 mAd541_1 mAd541_2 h3 j2 basic__key adr=541
Xkey@403 mAd520_1 mAd520_2 g3 j2 basic__key adr=520
Xkey@404 mAd657_1 mAd657_2 g5 j2 basic__key adr=657
Xkey@405 mAd636_1 mAd636_2 h5 j2 basic__key adr=636
Xkey@406 mAd762_1 mAd762_2 h7 Z10 basic__key adr=762
Xkey@407 mAd761_1 mAd761_2 g7 Z10 basic__key adr=761
Xkey@408 mAd750_1 mAd750_2 K13 Z10 basic__key adr=750
Xkey@409 mAd730_1 mAd730_2 K13 Z11 basic__key adr=730
Xkey@410 mAd741_1 mAd741_2 g7 Z11 basic__key adr=741
Xkey@411 mAd630_1 mAd630_2 K10 k3 basic__key adr=630
Xkey@412 mAd631_1 mAd631_2 K9 k3 basic__key adr=631
Xkey@413 mAd637_1 mAd637_2 g5 k2 basic__key adr=637
Xkey@414 mAd540_1 mAd540_2 g3 k2 basic__key adr=540
Xkey@415 mAd546_1 mAd546_2 K4 k1 basic__key adr=546
Xkey@416 mAd547_1 mAd547_2 K3 k1 basic__key adr=547
Xkey@417 mAd436_1 mAd436_2 g1 X11 basic__key adr=436
Xkey@418 mAd450_1 mAd450_2 K2 l1 basic__key adr=450
Xkey@419 mAd567_1 mAd567_2 K3 l1 basic__key adr=567
Xkey@420 mAd566_1 mAd566_2 K4 l1 basic__key adr=566
Xkey@421 mAd565_1 mAd565_2 K5 l1 basic__key adr=565
Xkey@422 mAd612_1 mAd612_2 K8 l3 basic__key adr=612
Xkey@423 mAd611_1 mAd611_2 K9 l3 basic__key adr=611
Xkey@424 mAd610_1 mAd610_2 K10 l3 basic__key adr=610
Xkey@425 mAd727_1 mAd727_2 K11 l3 basic__key adr=727
Xkey@426 mAd710_1 mAd710_2 K13 Z12 basic__key adr=710
Xkey@427 mAd700_1 mAd700_2 K13 X13 basic__key adr=700
Xkey@428 mAd711_1 mAd711_2 K12 X13 basic__key adr=711
Xkey@429 mAd717_1 mAd717_2 K11 X13 basic__key adr=717
Xkey@430 mAd600_1 mAd600_2 K10 X13 basic__key adr=600
Xkey@431 mAd601_1 mAd601_2 K9 X13 basic__key adr=601
Xkey@432 mAd602_1 mAd602_2 K8 X13 basic__key adr=602
Xkey@433 mAd607_1 mAd607_2 K7 X13 basic__key adr=607
Xkey@434 mAd570_1 mAd570_2 K6 X13 basic__key adr=570
Xkey@435 mAd575_1 mAd575_2 K5 X13 basic__key adr=575
Xkey@436 mAd576_1 mAd576_2 K4 X13 basic__key adr=576
Xkey@437 mAd577_1 mAd577_2 K3 X13 basic__key adr=577
Xkey@438 mAd460_1 mAd460_2 K2 X13 basic__key adr=460
Xkey@439 mAd466_1 mAd466_2 K1 X13 basic__key adr=466
.ENDS _5400TP094__CB

.global gnd

*** TOP LEVEL CELL: 123{sch}
.options filetype=ascii
.tran 0.1u 4u
.include "C:/IvanovFolder/PADIC/Spice64/models/soimod018.tec"
.global VDDA! VSSA!
.options method=gear reltol=0.01 itl4=500 altinit=10 RSHUNT=1.41G cshunt=1e-15 abstol=5u chgtol=2p vntol=5u trtol=7
XCB@1 CB@1_K0 CB@1_K1 CB@1_K10 CB@1_K11 CB@1_K12 CB@1_K13 CB@1_K2 CB@1_K3 CB@1_K4 CB@1_K5 CB@1_K6 CB@1_K7 CB@1_K8 CB@1_K9 CB@1_mAd000_1 CB@1_mAd000_2 CB@1_mAd001_1 CB@1_mAd001_2 CB@1_mAd002_1 CB@1_mAd002_2 CB@1_mAd003_1 CB@1_mAd003_2 CB@1_mAd004_1 CB@1_mAd004_2 CB@1_mAd005_1 CB@1_mAd005_2 CB@1_mAd006_1 CB@1_mAd006_2 CB@1_mAd007_1 CB@1_mAd007_2 CB@1_mAd010_1 CB@1_mAd010_2 CB@1_mAd011_1 CB@1_mAd011_2 CB@1_mAd012_1 CB@1_mAd012_2 CB@1_mAd013_1 CB@1_mAd013_2 CB@1_mAd014_1 CB@1_mAd014_2 CB@1_mAd015_1 
+CB@1_mAd015_2 CB@1_mAd016_1 CB@1_mAd016_2 CB@1_mAd017_1 CB@1_mAd017_2 CB@1_mAd020_1 CB@1_mAd020_2 CB@1_mAd021_1 CB@1_mAd021_2 CB@1_mAd022_1 CB@1_mAd022_2 CB@1_mAd023_1 CB@1_mAd023_2 CB@1_mAd024_1 CB@1_mAd024_2 CB@1_mAd025_1 CB@1_mAd025_2 CB@1_mAd026_1 CB@1_mAd026_2 CB@1_mAd027_1 CB@1_mAd027_2 CB@1_mAd030_1 CB@1_mAd030_2 CB@1_mAd031_1 CB@1_mAd031_2 CB@1_mAd032_1 CB@1_mAd032_2 CB@1_mAd033_1 CB@1_mAd033_2 CB@1_mAd034_1 CB@1_mAd034_2 CB@1_mAd035_1 CB@1_mAd035_2 CB@1_mAd036_1 CB@1_mAd036_2 CB@1_mAd037_1 
+CB@1_mAd037_2 CB@1_mAd040_1 CB@1_mAd040_2 CB@1_mAd041_1 CB@1_mAd041_2 CB@1_mAd042_1 CB@1_mAd042_2 CB@1_mAd043_1 CB@1_mAd043_2 CB@1_mAd044_1 CB@1_mAd044_2 CB@1_mAd045_1 CB@1_mAd045_2 CB@1_mAd046_1 CB@1_mAd046_2 CB@1_mAd047_1 CB@1_mAd047_2 CB@1_mAd050_1 CB@1_mAd050_2 CB@1_mAd051_1 CB@1_mAd051_2 CB@1_mAd052_1 CB@1_mAd052_2 CB@1_mAd053_1 CB@1_mAd053_2 CB@1_mAd054_1 CB@1_mAd054_2 CB@1_mAd055_1 CB@1_mAd055_2 CB@1_mAd056_1 CB@1_mAd056_2 CB@1_mAd057_1 CB@1_mAd057_2 CB@1_mAd060_1 CB@1_mAd060_2 CB@1_mAd066_1 
+CB@1_mAd066_2 CB@1_mAd067_1 CB@1_mAd067_2 CB@1_mAd100_1 CB@1_mAd100_2 CB@1_mAd101_1 CB@1_mAd101_2 CB@1_mAd102_1 CB@1_mAd102_2 CB@1_mAd110_1 CB@1_mAd110_2 CB@1_mAd111_1 CB@1_mAd111_2 CB@1_mAd112_1 CB@1_mAd112_2 CB@1_mAd113_1 CB@1_mAd113_2 CB@1_mAd114_1 CB@1_mAd114_2 CB@1_mAd115_1 CB@1_mAd115_2 CB@1_mAd116_1 CB@1_mAd116_2 CB@1_mAd117_1 CB@1_mAd117_2 CB@1_mAd120_1 CB@1_mAd120_2 CB@1_mAd121_1 CB@1_mAd121_2 CB@1_mAd122_1 CB@1_mAd122_2 CB@1_mAd123_1 CB@1_mAd123_2 CB@1_mAd124_1 CB@1_mAd124_2 CB@1_mAd125_1 
+CB@1_mAd125_2 CB@1_mAd126_1 CB@1_mAd126_2 CB@1_mAd127_1 CB@1_mAd127_2 CB@1_mAd130_1 CB@1_mAd130_2 CB@1_mAd131_1 CB@1_mAd131_2 CB@1_mAd132_1 CB@1_mAd132_2 CB@1_mAd133_1 CB@1_mAd133_2 CB@1_mAd134_1 CB@1_mAd134_2 CB@1_mAd135_1 CB@1_mAd135_2 CB@1_mAd136_1 CB@1_mAd136_2 CB@1_mAd137_1 CB@1_mAd137_2 CB@1_mAd140_1 CB@1_mAd140_2 CB@1_mAd141_1 CB@1_mAd141_2 CB@1_mAd142_1 CB@1_mAd142_2 CB@1_mAd143_1 CB@1_mAd143_2 CB@1_mAd144_1 CB@1_mAd144_2 CB@1_mAd145_1 CB@1_mAd145_2 CB@1_mAd146_1 CB@1_mAd146_2 CB@1_mAd147_1 
+CB@1_mAd147_2 CB@1_mAd150_1 CB@1_mAd150_2 CB@1_mAd151_1 CB@1_mAd151_2 CB@1_mAd152_1 CB@1_mAd152_2 CB@1_mAd153_1 CB@1_mAd153_2 CB@1_mAd154_1 CB@1_mAd154_2 CB@1_mAd155_1 CB@1_mAd155_2 CB@1_mAd156_1 CB@1_mAd156_2 CB@1_mAd157_1 CB@1_mAd157_2 CB@1_mAd160_1 CB@1_mAd160_2 CB@1_mAd161_1 CB@1_mAd161_2 CB@1_mAd162_1 CB@1_mAd162_2 CB@1_mAd163_1 CB@1_mAd163_2 CB@1_mAd164_1 CB@1_mAd164_2 CB@1_mAd165_1 CB@1_mAd165_2 CB@1_mAd166_1 CB@1_mAd166_2 CB@1_mAd167_1 CB@1_mAd167_2 CB@1_mAd170_1 CB@1_mAd170_2 CB@1_mAd171_1 
+CB@1_mAd171_2 CB@1_mAd172_1 CB@1_mAd172_2 CB@1_mAd173_1 CB@1_mAd173_2 CB@1_mAd175_1 CB@1_mAd175_2 CB@1_mAd176_1 CB@1_mAd176_2 CB@1_mAd177_1 CB@1_mAd177_2 CB@1_mAd200_1 CB@1_mAd200_2 CB@1_mAd201_1 CB@1_mAd201_2 CB@1_mAd202_1 CB@1_mAd202_2 CB@1_mAd204_1 CB@1_mAd204_2 CB@1_mAd205_1 CB@1_mAd205_2 CB@1_mAd206_1 CB@1_mAd206_2 CB@1_mAd207_1 CB@1_mAd207_2 CB@1_mAd210_1 CB@1_mAd210_2 CB@1_mAd211_1 CB@1_mAd211_2 CB@1_mAd212_1 CB@1_mAd212_2 CB@1_mAd213_1 CB@1_mAd213_2 CB@1_mAd214_1 CB@1_mAd214_2 CB@1_mAd215_1 
+CB@1_mAd215_2 CB@1_mAd216_1 CB@1_mAd216_2 CB@1_mAd217_1 CB@1_mAd217_2 CB@1_mAd220_1 CB@1_mAd220_2 CB@1_mAd221_1 CB@1_mAd221_2 CB@1_mAd222_1 CB@1_mAd222_2 CB@1_mAd223_1 CB@1_mAd223_2 CB@1_mAd224_1 CB@1_mAd224_2 CB@1_mAd225_1 CB@1_mAd225_2 CB@1_mAd226_1 CB@1_mAd226_2 CB@1_mAd227_1 CB@1_mAd227_2 CB@1_mAd230_1 CB@1_mAd230_2 CB@1_mAd231_1 CB@1_mAd231_2 CB@1_mAd232_1 CB@1_mAd232_2 CB@1_mAd233_1 CB@1_mAd233_2 CB@1_mAd234_1 CB@1_mAd234_2 CB@1_mAd235_1 CB@1_mAd235_2 CB@1_mAd236_1 CB@1_mAd236_2 CB@1_mAd237_1 
+CB@1_mAd237_2 CB@1_mAd240_1 CB@1_mAd240_2 CB@1_mAd241_1 CB@1_mAd241_2 CB@1_mAd242_1 CB@1_mAd242_2 CB@1_mAd243_1 CB@1_mAd243_2 CB@1_mAd244_1 CB@1_mAd244_2 CB@1_mAd245_1 CB@1_mAd245_2 CB@1_mAd246_1 CB@1_mAd246_2 CB@1_mAd247_1 CB@1_mAd247_2 CB@1_mAd250_1 CB@1_mAd250_2 CB@1_mAd251_1 CB@1_mAd251_2 CB@1_mAd252_1 CB@1_mAd252_2 CB@1_mAd253_1 CB@1_mAd253_2 CB@1_mAd254_1 CB@1_mAd254_2 CB@1_mAd255_1 CB@1_mAd255_2 CB@1_mAd256_1 CB@1_mAd256_2 CB@1_mAd257_1 CB@1_mAd257_2 CB@1_mAd260_1 CB@1_mAd260_2 CB@1_mAd261_1 
+CB@1_mAd261_2 CB@1_mAd262_1 CB@1_mAd262_2 CB@1_mAd263_1 CB@1_mAd263_2 CB@1_mAd264_1 CB@1_mAd264_2 CB@1_mAd265_1 CB@1_mAd265_2 CB@1_mAd266_1 CB@1_mAd266_2 CB@1_mAd267_1 CB@1_mAd267_2 CB@1_mAd275_1 CB@1_mAd275_2 CB@1_mAd276_1 CB@1_mAd276_2 CB@1_mAd277_1 CB@1_mAd277_2 CB@1_mAd300_1 CB@1_mAd300_2 CB@1_mAd310_1 CB@1_mAd310_2 CB@1_mAd311_1 CB@1_mAd311_2 CB@1_mAd317_1 CB@1_mAd317_2 CB@1_mAd320_1 CB@1_mAd320_2 CB@1_mAd321_1 CB@1_mAd321_2 CB@1_mAd322_1 CB@1_mAd322_2 CB@1_mAd323_1 CB@1_mAd323_2 CB@1_mAd324_1 
+CB@1_mAd324_2 CB@1_mAd325_1 CB@1_mAd325_2 CB@1_mAd326_1 CB@1_mAd326_2 CB@1_mAd327_1 CB@1_mAd327_2 CB@1_mAd330_1 CB@1_mAd330_2 CB@1_mAd331_1 CB@1_mAd331_2 CB@1_mAd332_1 CB@1_mAd332_2 CB@1_mAd333_1 CB@1_mAd333_2 CB@1_mAd334_1 CB@1_mAd334_2 CB@1_mAd335_1 CB@1_mAd335_2 CB@1_mAd336_1 CB@1_mAd336_2 CB@1_mAd337_1 CB@1_mAd337_2 CB@1_mAd340_1 CB@1_mAd340_2 CB@1_mAd341_1 CB@1_mAd341_2 CB@1_mAd342_1 CB@1_mAd342_2 CB@1_mAd343_1 CB@1_mAd343_2 CB@1_mAd344_1 CB@1_mAd344_2 CB@1_mAd345_1 CB@1_mAd345_2 CB@1_mAd346_1 
+CB@1_mAd346_2 CB@1_mAd347_1 CB@1_mAd347_2 CB@1_mAd350_1 CB@1_mAd350_2 CB@1_mAd351_1 CB@1_mAd351_2 CB@1_mAd352_1 CB@1_mAd352_2 CB@1_mAd353_1 CB@1_mAd353_2 CB@1_mAd354_1 CB@1_mAd354_2 CB@1_mAd355_1 CB@1_mAd355_2 CB@1_mAd356_1 CB@1_mAd356_2 CB@1_mAd357_1 CB@1_mAd357_2 CB@1_mAd360_1 CB@1_mAd360_2 CB@1_mAd361_1 CB@1_mAd361_2 CB@1_mAd362_1 CB@1_mAd362_2 CB@1_mAd363_1 CB@1_mAd363_2 CB@1_mAd364_1 CB@1_mAd364_2 CB@1_mAd365_1 CB@1_mAd365_2 CB@1_mAd366_1 CB@1_mAd366_2 CB@1_mAd367_1 CB@1_mAd367_2 CB@1_mAd371_1 
+CB@1_mAd371_2 CB@1_mAd372_1 CB@1_mAd372_2 CB@1_mAd373_1 CB@1_mAd373_2 CB@1_mAd374_1 CB@1_mAd374_2 CB@1_mAd375_1 CB@1_mAd375_2 CB@1_mAd376_1 CB@1_mAd376_2 CB@1_mAd377_1 CB@1_mAd377_2 CB@1_mAd400_1 CB@1_mAd400_2 CB@1_mAd401_1 CB@1_mAd401_2 CB@1_mAd402_1 CB@1_mAd402_2 CB@1_mAd403_1 CB@1_mAd403_2 CB@1_mAd404_1 CB@1_mAd404_2 CB@1_mAd405_1 CB@1_mAd405_2 CB@1_mAd406_1 CB@1_mAd406_2 CB@1_mAd407_1 CB@1_mAd407_2 CB@1_mAd410_1 CB@1_mAd410_2 CB@1_mAd411_1 CB@1_mAd411_2 CB@1_mAd412_1 CB@1_mAd412_2 CB@1_mAd413_1 
+CB@1_mAd413_2 CB@1_mAd414_1 CB@1_mAd414_2 CB@1_mAd415_1 CB@1_mAd415_2 CB@1_mAd416_1 CB@1_mAd416_2 CB@1_mAd417_1 CB@1_mAd417_2 CB@1_mAd420_1 CB@1_mAd420_2 CB@1_mAd421_1 CB@1_mAd421_2 CB@1_mAd422_1 CB@1_mAd422_2 CB@1_mAd423_1 CB@1_mAd423_2 CB@1_mAd424_1 CB@1_mAd424_2 CB@1_mAd425_1 CB@1_mAd425_2 CB@1_mAd426_1 CB@1_mAd426_2 CB@1_mAd427_1 CB@1_mAd427_2 CB@1_mAd430_1 CB@1_mAd430_2 CB@1_mAd431_1 CB@1_mAd431_2 CB@1_mAd432_1 CB@1_mAd432_2 CB@1_mAd433_1 CB@1_mAd433_2 CB@1_mAd434_1 CB@1_mAd434_2 CB@1_mAd435_1 
+CB@1_mAd435_2 CB@1_mAd436_1 CB@1_mAd436_2 CB@1_mAd437_1 CB@1_mAd437_2 CB@1_mAd440_1 CB@1_mAd440_2 CB@1_mAd441_1 CB@1_mAd441_2 CB@1_mAd442_1 CB@1_mAd442_2 CB@1_mAd443_1 CB@1_mAd443_2 CB@1_mAd444_1 CB@1_mAd444_2 CB@1_mAd445_1 CB@1_mAd445_2 CB@1_mAd446_1 CB@1_mAd446_2 CB@1_mAd447_1 CB@1_mAd447_2 CB@1_mAd450_1 CB@1_mAd450_2 CB@1_mAd451_1 CB@1_mAd451_2 CB@1_mAd452_1 CB@1_mAd452_2 CB@1_mAd453_1 CB@1_mAd453_2 CB@1_mAd454_1 CB@1_mAd454_2 CB@1_mAd455_1 CB@1_mAd455_2 CB@1_mAd456_1 CB@1_mAd456_2 CB@1_mAd457_1 
+CB@1_mAd457_2 CB@1_mAd460_1 CB@1_mAd460_2 CB@1_mAd466_1 CB@1_mAd466_2 CB@1_mAd467_1 CB@1_mAd467_2 CB@1_mAd500_1 CB@1_mAd500_2 CB@1_mAd501_1 CB@1_mAd501_2 CB@1_mAd502_1 CB@1_mAd502_2 CB@1_mAd508_1 CB@1_mAd508_2 CB@1_mAd509_1 CB@1_mAd509_2 CB@1_mAd512_1 CB@1_mAd512_2 CB@1_mAd513_1 CB@1_mAd513_2 CB@1_mAd514_1 CB@1_mAd514_2 CB@1_mAd515_1 CB@1_mAd515_2 CB@1_mAd516_1 CB@1_mAd516_2 CB@1_mAd517_1 CB@1_mAd517_2 CB@1_mAd520_1 CB@1_mAd520_2 CB@1_mAd521_1 CB@1_mAd521_2 CB@1_mAd522_1 CB@1_mAd522_2 CB@1_mAd523_1 
+CB@1_mAd523_2 CB@1_mAd524_1 CB@1_mAd524_2 CB@1_mAd525_1 CB@1_mAd525_2 CB@1_mAd526_1 CB@1_mAd526_2 CB@1_mAd527_1 CB@1_mAd527_2 CB@1_mAd530_1 CB@1_mAd530_2 CB@1_mAd531_1 CB@1_mAd531_2 CB@1_mAd532_1 CB@1_mAd532_2 CB@1_mAd533_1 CB@1_mAd533_2 CB@1_mAd534_1 CB@1_mAd534_2 CB@1_mAd535_1 CB@1_mAd535_2 CB@1_mAd536_1 CB@1_mAd536_2 CB@1_mAd537_1 CB@1_mAd537_2 CB@1_mAd540_1 CB@1_mAd540_2 CB@1_mAd541_1 CB@1_mAd541_2 CB@1_mAd542_1 CB@1_mAd542_2 CB@1_mAd543_1 CB@1_mAd543_2 CB@1_mAd544_1 CB@1_mAd544_2 CB@1_mAd545_1 
+CB@1_mAd545_2 CB@1_mAd546_1 CB@1_mAd546_2 CB@1_mAd547_1 CB@1_mAd547_2 CB@1_mAd550_1 CB@1_mAd550_2 CB@1_mAd551_1 CB@1_mAd551_2 CB@1_mAd552_1 CB@1_mAd552_2 CB@1_mAd553_1 CB@1_mAd553_2 CB@1_mAd554_1 CB@1_mAd554_2 CB@1_mAd555_1 CB@1_mAd555_2 CB@1_mAd556_1 CB@1_mAd556_2 CB@1_mAd557_1 CB@1_mAd557_2 CB@1_mAd560_1 CB@1_mAd560_2 CB@1_mAd561_1 CB@1_mAd561_2 CB@1_mAd562_1 CB@1_mAd562_2 CB@1_mAd563_1 CB@1_mAd563_2 CB@1_mAd564_1 CB@1_mAd564_2 CB@1_mAd565_1 CB@1_mAd565_2 CB@1_mAd566_1 CB@1_mAd566_2 CB@1_mAd567_1 
+CB@1_mAd567_2 CB@1_mAd570_1 CB@1_mAd570_2 CB@1_mAd571_1 CB@1_mAd571_2 CB@1_mAd572_1 CB@1_mAd572_2 CB@1_mAd573_1 CB@1_mAd573_2 CB@1_mAd575_1 CB@1_mAd575_2 CB@1_mAd576_1 CB@1_mAd576_2 CB@1_mAd577_1 CB@1_mAd577_2 CB@1_mAd600_1 CB@1_mAd600_2 CB@1_mAd601_1 CB@1_mAd601_2 CB@1_mAd602_1 CB@1_mAd602_2 CB@1_mAd604_1 CB@1_mAd604_2 CB@1_mAd605_1 CB@1_mAd605_2 CB@1_mAd606_1 CB@1_mAd606_2 CB@1_mAd607_1 CB@1_mAd607_2 CB@1_mAd610_1 CB@1_mAd610_2 CB@1_mAd611_1 CB@1_mAd611_2 CB@1_mAd612_1 CB@1_mAd612_2 CB@1_mAd613_1 
+CB@1_mAd613_2 CB@1_mAd614_1 CB@1_mAd614_2 CB@1_mAd615_1 CB@1_mAd615_2 CB@1_mAd616_1 CB@1_mAd616_2 CB@1_mAd617_1 CB@1_mAd617_2 CB@1_mAd620_1 CB@1_mAd620_2 CB@1_mAd621_1 CB@1_mAd621_2 CB@1_mAd622_1 CB@1_mAd622_2 CB@1_mAd623_1 CB@1_mAd623_2 CB@1_mAd624_1 CB@1_mAd624_2 CB@1_mAd625_1 CB@1_mAd625_2 CB@1_mAd626_1 CB@1_mAd626_2 CB@1_mAd627_1 CB@1_mAd627_2 CB@1_mAd630_1 CB@1_mAd630_2 CB@1_mAd631_1 CB@1_mAd631_2 CB@1_mAd632_1 CB@1_mAd632_2 CB@1_mAd633_1 CB@1_mAd633_2 CB@1_mAd634_1 CB@1_mAd634_2 CB@1_mAd635_1 
+CB@1_mAd635_2 CB@1_mAd636_1 CB@1_mAd636_2 CB@1_mAd637_1 CB@1_mAd637_2 CB@1_mAd640_1 CB@1_mAd640_2 CB@1_mAd641_1 CB@1_mAd641_2 CB@1_mAd642_1 CB@1_mAd642_2 CB@1_mAd643_1 CB@1_mAd643_2 CB@1_mAd644_1 CB@1_mAd644_2 CB@1_mAd645_1 CB@1_mAd645_2 CB@1_mAd646_1 CB@1_mAd646_2 CB@1_mAd647_1 CB@1_mAd647_2 CB@1_mAd650_1 CB@1_mAd650_2 CB@1_mAd651_1 CB@1_mAd651_2 CB@1_mAd652_1 CB@1_mAd652_2 CB@1_mAd653_1 CB@1_mAd653_2 CB@1_mAd654_1 CB@1_mAd654_2 CB@1_mAd655_1 CB@1_mAd655_2 CB@1_mAd656_1 CB@1_mAd656_2 CB@1_mAd657_1 
+CB@1_mAd657_2 CB@1_mAd660_1 CB@1_mAd660_2 CB@1_mAd661_1 CB@1_mAd661_2 CB@1_mAd662_1 CB@1_mAd662_2 CB@1_mAd663_1 CB@1_mAd663_2 CB@1_mAd664_1 CB@1_mAd664_2 CB@1_mAd665_1 CB@1_mAd665_2 CB@1_mAd666_1 CB@1_mAd666_2 CB@1_mAd667_1 CB@1_mAd667_2 CB@1_mAd675_1 CB@1_mAd675_2 CB@1_mAd676_1 CB@1_mAd676_2 CB@1_mAd677_1 CB@1_mAd677_2 CB@1_mAd700_1 CB@1_mAd700_2 CB@1_mAd710_1 CB@1_mAd710_2 CB@1_mAd711_1 CB@1_mAd711_2 CB@1_mAd717_1 CB@1_mAd717_2 CB@1_mAd720_1 CB@1_mAd720_2 CB@1_mAd721_1 CB@1_mAd721_2 CB@1_mAd722_1 
+CB@1_mAd722_2 CB@1_mAd723_1 CB@1_mAd723_2 CB@1_mAd724_1 CB@1_mAd724_2 CB@1_mAd725_1 CB@1_mAd725_2 CB@1_mAd726_1 CB@1_mAd726_2 CB@1_mAd727_1 CB@1_mAd727_2 CB@1_mAd730_1 CB@1_mAd730_2 CB@1_mAd731_1 CB@1_mAd731_2 CB@1_mAd732_1 CB@1_mAd732_2 CB@1_mAd733_1 CB@1_mAd733_2 CB@1_mAd734_1 CB@1_mAd734_2 CB@1_mAd735_1 CB@1_mAd735_2 CB@1_mAd736_1 CB@1_mAd736_2 CB@1_mAd737_1 CB@1_mAd737_2 CB@1_mAd740_1 CB@1_mAd740_2 CB@1_mAd741_1 CB@1_mAd741_2 CB@1_mAd742_1 CB@1_mAd742_2 CB@1_mAd743_1 CB@1_mAd743_2 CB@1_mAd744_1 
+CB@1_mAd744_2 CB@1_mAd745_1 CB@1_mAd745_2 CB@1_mAd746_1 CB@1_mAd746_2 CB@1_mAd747_1 CB@1_mAd747_2 CB@1_mAd750_1 CB@1_mAd750_2 CB@1_mAd751_1 CB@1_mAd751_2 CB@1_mAd752_1 CB@1_mAd752_2 CB@1_mAd753_1 CB@1_mAd753_2 CB@1_mAd754_1 CB@1_mAd754_2 CB@1_mAd755_1 CB@1_mAd755_2 CB@1_mAd756_1 CB@1_mAd756_2 CB@1_mAd757_1 CB@1_mAd757_2 CB@1_mAd760_1 CB@1_mAd760_2 CB@1_mAd761_1 CB@1_mAd761_2 CB@1_mAd762_1 CB@1_mAd762_2 CB@1_mAd763_1 CB@1_mAd763_2 CB@1_mAd764_1 CB@1_mAd764_2 CB@1_mAd765_1 CB@1_mAd765_2 CB@1_mAd766_1 
+CB@1_mAd766_2 CB@1_mAd767_1 CB@1_mAd767_2 CB@1_mAd771_1 CB@1_mAd771_2 CB@1_mAd772_1 CB@1_mAd772_2 CB@1_mAd773_1 CB@1_mAd773_2 CB@1_mAd774_1 CB@1_mAd774_2 CB@1_mAd775_1 CB@1_mAd775_2 CB@1_mAd776_1 CB@1_mAd776_2 CB@1_mAd777_1 CB@1_mAd777_2 CB@1_X0 CB@1_X1 CB@1_X10 CB@1_X11 CB@1_X12 CB@1_X13 CB@1_X2 CB@1_X3 CB@1_X4 CB@1_X5 CB@1_X6 CB@1_X7 CB@1_X8 CB@1_X9 CB@1_Y1 CB@1_Y10 CB@1_Y11 CB@1_Y12 CB@1_Y2 CB@1_Y3 CB@1_Y4 CB@1_Y5 CB@1_Y6 CB@1_Y7 CB@1_Y8 CB@1_Y9 CB@1_Z1 CB@1_Z10 CB@1_Z11 CB@1_Z12 CB@1_Z2 CB@1_Z3 CB@1_Z4 
+CB@1_Z5 CB@1_Z6 CB@1_Z7 CB@1_Z8 CB@1_Z9 _5400TP094__CB
.END
